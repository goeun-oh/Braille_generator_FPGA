/*******************************************************************************
Author: joohan.kim (https://blog.naver.com/chacagea)
Associated Filename: cnn_core.v
Purpose: verilog code to understand the CNN operation
License : https://github.com/matbi86/matbi_fpga_season_1/blob/main/LICENSE
Revision History: February 13, 2020 - initial release
*******************************************************************************/

`include "timescale.v"
`include "defines_cnn_core.v"

module cnn_kernel (
    // Clock & Reset
input                               	clk         	,
input                               	reset_n     	,

//5x5x7
input     [`KX*`KY*`W_BW-1 : 0] 	    i_cnn_weight 	,
input                                   i_in_valid  	,
input     [`KX*`KY*`ST2_Conv_IBW-1 : 0] i_in_fmap    	,
output                                  o_ot_valid  	,
output    [`AK_BW-1 : 0]  			    o_ot_kernel_acc           
    );

localparam LATENCY = 2;




//==============================================================================
// Data Enable Signals 
//==============================================================================
wire    [LATENCY-1 : 0] 	ce;
reg     [LATENCY-1 : 0] 	r_valid;
always @(posedge clk or negedge reset_n) begin
    if(!reset_n) begin
        r_valid   <= {LATENCY{1'b0}};
    end else begin
        r_valid[LATENCY-2]  <= i_in_valid;
        r_valid[LATENCY-1]  <= r_valid[LATENCY-2];
    end
end

assign	ce = r_valid;

//==============================================================================
// mul = fmap * weight
//==============================================================================

wire      [`KY*`KX*`M_BW-1 : 0]    mul  ;
reg       [`KY*`KX*`M_BW-1 : 0]    r_mul;

genvar mul_idx;
generate
	//커널사이즈(5x5만큼 한번의 곱셈하기 위함)
	for(mul_idx = 0; mul_idx < `KY*`KX; mul_idx = mul_idx + 1) begin : gen_mul
		assign  mul[mul_idx * `M_BW +: `M_BW]	= i_in_fmap[mul_idx * `ST2_Conv_IBW +: `ST2_Conv_IBW] * i_cnn_weight[mul_idx * `W_BW +: `W_BW];
	
		always @(posedge clk or negedge reset_n) begin
		    if(!reset_n) begin
		        r_mul[mul_idx * `M_BW +: `M_BW] <= {`M_BW{1'b0}};
		    end else if(i_in_valid)begin
		        r_mul[mul_idx * `M_BW +: `M_BW] <= mul[mul_idx * `M_BW +: `M_BW];
		    end
		end
	end
endgenerate

reg       [`AK_BW-1 : 0]    acc_kernel 	;
reg       [`AK_BW-1 : 0]    r_acc_kernel   ;

integer acc_idx;
generate
	always @ (*) begin
		acc_kernel[0 +: `AK_BW]= {`AK_BW{1'b0}};
		for(acc_idx =0; acc_idx < `KY*`KX; acc_idx = acc_idx +1) begin
			acc_kernel[0 +: `AK_BW] = acc_kernel[0 +: `AK_BW] + r_mul[acc_idx*`M_BW +: `M_BW]; 
		end
	end
	always @(posedge clk or negedge reset_n) begin
	    if(!reset_n) begin
	        r_acc_kernel[0 +: `AK_BW] <= {`AK_BW{1'b0}};
	    end else if(ce[LATENCY-2])begin
	        r_acc_kernel[0 +: `AK_BW] <= acc_kernel[0 +: `AK_BW];
	    end
	end
endgenerate

assign o_ot_valid = r_valid[LATENCY-1];
assign o_ot_kernel_acc = r_acc_kernel;

endmodule
