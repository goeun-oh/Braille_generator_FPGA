`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2025/07/20 07:17:32
// Design Name: 
// Module Name: conv2_weight_rom
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

`include "defines_cnn_core.v"


module conv2_weight_rom #(
    parameter CHANNEL_ID = 0
)(
    output reg signed [`ST2_Conv_CO * `KX * `KY * `W_BW-1:0] weight   //3x3x5x5x(7bit) 중 1개를 3x5x5x(7bit)로 출력
);

initial begin
     case (CHANNEL_ID)
        0: begin
                weight = {
                    7'd33, 7'd9, 7'd9, -7'd7, 7'd0,
                    7'd29, 7'd22, -7'd13, 7'd26, 7'd34,
                    7'd15, 7'd5, 7'd26, 7'd37, 7'd46,
                    7'd19, 7'd27, 7'd31, 7'd37, 7'd33,
                    -7'd2, 7'd11, 7'd7, -7'd5, -7'd3,

                    7'd14, 7'd16, 7'd14, 7'd17, 7'd34,
                    7'd15, -7'd5, 7'd15, 7'd26, 7'd15,
                    -7'd31, 7'd13, -7'd1, 7'd1, 7'd17,
                    -7'd19, -7'd9, -7'd24, -7'd15, -7'd2,
                    -7'd29, -7'd31, -7'd5, -7'd22, -7'd17,

                    7'd4, -7'd17, 7'd4, -7'd7, -7'd7,
                    7'd35, -7'd27, -7'd36, -7'd16, 7'd25,
                    7'd30, 7'd27, 7'd14, 7'd39, 7'd44,
                    7'd47, 7'd41, 7'd45, 7'd37, 7'd31,
                    7'd46, 7'd52, 7'd27, -7'd4, -7'd5
                };
            end
        1: begin
                weight = {
                    -7'd16, -7'd29, -7'd37, -7'd6, -7'd24,
                    -7'd27, -7'd27, -7'd2, 7'd4, 7'd5,
                    -7'd9, -7'd4, -7'd1, -7'd7, 7'd17,
                    7'd11, 7'd7, -7'd20, -7'd6, 7'd4,
                    7'd25, 7'd7, 7'd15, -7'd5, 7'd16,

                    -7'd1, -7'd30, -7'd10, 7'd22, 7'd10,
                    7'd13, 7'd11, -7'd6, 7'd1, 7'd37,
                    7'd34, 7'd12, 7'd6, 7'd7, 7'd30,
                    7'd33, 7'd26, 7'd30, 7'd9, 7'd23,
                    7'd51, 7'd25, 7'd29, 7'd16, 7'd9,

                    -7'd27, 7'd6, -7'd7, -7'd20, -7'd53,
                    -7'd34, -7'd20, 7'd3, -7'd4, -7'd47,
                    -7'd45, -7'd40, -7'd7, 7'd6, 7'd5,
                    -7'd66, -7'd56, -7'd52, -7'd35, -7'd27,
                    -7'd41, -7'd45, -7'd41, -7'd47, -7'd11
                };
            end
        2: begin
                weight = {
                    -7'd9, 7'd5, 7'd7, 7'd13, -7'd10,
                    -7'd7, -7'd16, -7'd2, 7'd10, 7'd3,
                    -7'd4, 7'd11, 7'd3, -7'd12, 7'd7,
                    7'd1, -7'd13, 7'd1, 7'd1, -7'd1,
                    -7'd10, -7'd14, -7'd15, 7'd0, -7'd6,

                    7'd11, 7'd11, -7'd7, -7'd13, 7'd4,
                    -7'd15, 7'd6, -7'd15, -7'd9, 7'd6,
                    -7'd9, -7'd7, 7'd0, -7'd1, -7'd10,
                    -7'd9, 7'd3, 7'd1, 7'd2, -7'd9,
                    -7'd2, -7'd4, -7'd3, 7'd2, -7'd15,

                    7'd5, 7'd2, 7'd3, -7'd15, -7'd9,
                    -7'd13, 7'd2, 7'd2, -7'd7, -7'd9,
                    7'd1, 7'd7, -7'd4, -7'd1, -7'd15,
                    7'd10, -7'd3, 7'd11, -7'd13, 7'd10,
                    -7'd7, 7'd1, 7'd9, -7'd12, -7'd5
                };
            end
        endcase
end


endmodule
