`timescale 1ns / 1ps
module display_lev1 (

    output logic [3:0] test_led,

    input logic pclk,  // 25MHz
    input logic reset,
    // VGA Controller side
    input logic [9:0] x_pixel,
    input logic [9:0] y_pixel,
    input logic [3:0] cam_r,  // 카메라 red 포트
    input logic [3:0] cam_g,  // 카메라 green 포트
    input logic [3:0] cam_b,  // 카메라 blue 포트
    // export side
    output logic slave_done,        // 한 라운드의 게임이 끝나면 알려주는 신호호
    output logic [3:0] red_port,  // vga red 포트
    output logic [3:0] green_port,  // vga green 포트
    output logic [3:0] blue_port,  // vga blue 포트

    // Control Board side
    input logic sw,  // start 신호 + 레벨 알려줄때 done 신호
    input logic [1:0] lvl,  // level 1,2,3
    input logic [7:0] question,  // 게임 RGB 값 받는 신호, 3가지 색깔 4개
    input logic give_done,

    // Color Detect side
    output logic countdown_done,    // 카운트다운이 7->0 되면 알려주는 신호

    // Color Comparison side
    input  logic comparison_done,
    output logic give_comparison_done,
    input  logic [1:0] win_lose,   // 게임 맞혔다 틀렸다 신호 , win_lose초기화 상태는 0으로 해주세요!!!

    // piezo
    output logic [1:0] startcount,
    output logic [3:0] countdown,
    output logic bgm_enable // IDLE bgm

);
  logic [63:0] Wout_bitmap [0:63] = {
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000111111111110000000000001111111111100000000000011111111111000,
    64'b0001111111111111000000000011111111111110000000000111111111111100,
    64'b0001111111111111000000000111111111111111000000001111111111111110,
    64'b0011111000001111100000001111110000011111000000001111100000111110,
    64'b0111110000000111110000001111100000001111100000011111000000011111,
    64'b0111110000000111110000001111000000000111100000011110000000001111,
    64'b0111100000000011110000001110000000000111110000011110000000001111,
    64'b0111000011100001110000011110001111000011110000111100001110000111,
    64'b0111000011100001111000011110001111100011110000111100011111000111,
    64'b0111000111110001111000111110001111100001110000111100011111000111,
    64'b0111000111110001111000111100011111110001111000111000011111000111,
    64'b0111000111111000111000111100011111110001111001111000111111000111,
    64'b0111000111111000111100111000011111110001111101111000111111000111,
    64'b0111000011111000111101111000011101111000111101111001111111001111,
    64'b0111100011111000111111111000111101111000111101110001111110001111,
    64'b0111100011111100011111111000111101111000011111110001111110001111,
    64'b0111100011111100011111110001111111111000011111110001111100001110,
    64'b0011110001111110001111110001111111111100011111110001111100001110,
    64'b0011110001111110001111110001111111111100011111100011111100011110,
    64'b0011110000111110001111100011111101111110001111000111111000111110,
    64'b0001111000111111001111100011111101111110001111000111111000111110,
    64'b0001111000111111000111100011111100111110001111000111110000111100,
    64'b0001111100011111000111000111111000111110001111000111110000111000,
    64'b0000111100011111000011000111111000111111000111001111110001111000,
    64'b0000111100011111000011000111110000111111000110001111110001111000,
    64'b0000011100011111100011000111110000011111100010001111100011111000,
    64'b0000011110001111100010001111110000011111100000001111100011110000,
    64'b0000011110001111110000001111110000011111100000001111100011110000,
    64'b0000011111000111110000011111100000011111100000011111100011100000,
    64'b0000001111000111110000011111100010001111110000011111000111100000,
    64'b0000001111000111110000011111100010001111110000111111000111100000,
    64'b0000000111000111111000011111100011000111110000111110001111100000,
    64'b0000000111100111111000011111000111000111110000111110001111000000,
    64'b0000000111100011111100111111000111000111110000111110001111000000,
    64'b0000000111100011111100111110001111000111111000111110001110000000,
    64'b0000000011100001111100111110001111100011111101111100011110000000,
    64'b0000000011110001111101111110001111100001111111111000011110000000,
    64'b0000000011110001111111111100011111100001111111111000011110000000,
    64'b0000000011111000111111111100011111110001111111111000011100000000,
    64'b0000000001111000111111111000011111110001111101111000111100000000,
    64'b0000000001111000111101111000011111111000111101111001111100000000,
    64'b0000000000111000111111111000111101111000111101110001111100000000,
    64'b0000000000111100011111111000111101111000011111110001111000000000,
    64'b0000000000111100011111110001111100111000011111110001110000000000,
    64'b0000000000111110001111110001111000111000011111110001110000000000,
    64'b0000000000011110001111100001111000111100011111100011110000000000,
    64'b0000000000011110001111100001110000111100001111000011110000000000,
    64'b0000000000001110000011000011110000111110001111000111110000000000,
    64'b0000000000001111000000000011110000011110000000000111100000000000,
    64'b0000000000001111000000000111110000011110000000000111100000000000,
    64'b0000000000001111100000000111100000001111000000001111000000000000,
    64'b0000000000000111111111111111100000001111111111111111000000000000,
    64'b0000000000000111111111111111000000001111111111111111000000000000,
    64'b0000000000000011111111111111000000000111111111111110000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000
};

logic [63:0] Wmid_bitmap [0:63] = {
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000111110000000000000000001111100000000000000000011111000000,
    64'b0000001111111000000000000000011111110000000000000000111111100000,
    64'b0000001111111000000000000000111111111000000000000001111111110000,
    64'b0000011111111100000000000001111111111000000000000001111111110000,
    64'b0000111100011110000000000001110000111100000000000011110001111000,
    64'b0000111100011110000000000001110000011100000000000011100000111000,
    64'b0000111000001110000000000001110000011110000000000011100000111000,
    64'b0000111000001110000000000011100000001110000000000111100000111000,
    64'b0000111000000111000000000011100000001110000000000111000000111000,
    64'b0000111000000111000000000111100000001110000000000111000000111000,
    64'b0000111100000111000000000111100000000111000000000110000000110000,
    64'b0000011100000111000000000111000000000111000000001110000001110000,
    64'b0000011100000011100000000111000000000111100000001110000001110000,
    64'b0000011100000011100000001110000000000111100000001110000011110000,
    64'b0000001110000001110000001110000000000011100000001110000011110000,
    64'b0000001110000001110000001110000000000011100000011100000011100000,
    64'b0000001111000001110000011100000010000001110000111000000111000000,
    64'b0000000111000000110000011100000010000001110000111000000111000000,
    64'b0000000111000000111000011100000011000001110000111000001111000000,
    64'b0000000011100000111000111000000111000001110000111000001111000000,
    64'b0000000011100000111100111000000111000000111000110000001110000000,
    64'b0000000011100000111100111000001111000000111001110000001110000000,
    64'b0000000011100000011100111000001111100000011101110000011100000000,
    64'b0000000001110000011101110000001111100000011111110000011100000000,
    64'b0000000001110000001111110000001111100000011111110000011100000000,
    64'b0000000000111000001111100000011111100000011111100000011100000000,
    64'b0000000000111000001111100000011101110000001111100000111000000000,
    64'b0000000000111000001111100000011101110000001111000000111000000000,
    64'b0000000000111000000111100000011100111000001111000001110000000000,
    64'b0000000000011000000111100000111000111000001111000001110000000000,
    64'b0000000000011100000011000000111000111000001111000001110000000000,
    64'b0000000000011100000011000001110000111000000111000001110000000000,
    64'b0000000000011110000011000001110000011100000010000011100000000000,
    64'b0000000000001110000010000001110000011110000000000111100000000000,
    64'b0000000000001110000000000011100000011110000000000111100000000000,
    64'b0000000000000111000000000011100000001110000000000111100000000000,
    64'b0000000000000111000000000111100000001110000000000111000000000000,
    64'b0000000000000111000000000111100000000111000000000110000000000000,
    64'b0000000000000111000000000111000000000111000000001110000000000000,
    64'b0000000000000011100000000111000000000111100000001110000000000000,
    64'b0000000000000011100000001110000000000111100000001110000000000000,
    64'b0000000000000001110000001110000000000111100000001110000000000000,
    64'b0000000000000001110000011110000000000011100000011100000000000000,
    64'b0000000000000001110000011110000000000011110000111100000000000000,
    64'b0000000000000001111100111100000000000001110000111000000000000000,
    64'b0000000000000000111111111100000000000001111111111000000000000000,
    64'b0000000000000000111111111000000000000001111111111000000000000000,
    64'b0000000000000000011111111000000000000000111111110000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000
};

logic [63:0] Win_bitmap [0:63] = {
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000011100000000000000000001111000000000000000000001110000000,
    64'b0000000011100000000000000000001111100000000000000000011111000000,
    64'b0000000111110000000000000000001111100000000000000000011111000000,
    64'b0000000111110000000000000000011111110000000000000000011111000000,
    64'b0000000111111000000000000000011111110000000000000000111111000000,
    64'b0000000111111000000000000000011111110000000000000000111111000000,
    64'b0000000011111000000000000000011111111000000000000001111111000000,
    64'b0000000011111000000000000000111111111000000000000001111110000000,
    64'b0000000011111100000000000000111111111000000000000001111110000000,
    64'b0000000011111100000000000001111111111000000000000001111100000000,
    64'b0000000001111110000000000001111111111100000000000001111100000000,
    64'b0000000001111110000000000001111111111100000000000011111100000000,
    64'b0000000000111110000000000011111101111110000000000111111000000000,
    64'b0000000000111111000000000011111101111110000000000111111000000000,
    64'b0000000000111111000000000011111100111110000000000111110000000000,
    64'b0000000000011111000000000111111000111110000000000111110000000000,
    64'b0000000000011111000000000111111000111111000000001111110000000000,
    64'b0000000000011111000000000111110000111111000000001111110000000000,
    64'b0000000000011111100000000111110000011111100000001111100000000000,
    64'b0000000000001111100000001111110000011111100000001111100000000000,
    64'b0000000000001111110000001111110000011111100000001111100000000000,
    64'b0000000000000111110000011111100000011111100000011111100000000000,
    64'b0000000000000111110000011111100000001111110000011111000000000000,
    64'b0000000000000111110000011111100000001111110000111111000000000000,
    64'b0000000000000111111000011111100000000111110000111110000000000000,
    64'b0000000000000111111000011111000000000111110000111110000000000000,
    64'b0000000000000011111100111111000000000111110000111110000000000000,
    64'b0000000000000011111100111110000000000111111000111110000000000000,
    64'b0000000000000001111100111110000000000011111101111100000000000000,
    64'b0000000000000001111101111110000000000001111111111000000000000000,
    64'b0000000000000001111111111100000000000001111111111000000000000000,
    64'b0000000000000000111111111100000000000001111111111000000000000000,
    64'b0000000000000000111111111000000000000001111111111000000000000000,
    64'b0000000000000000111111111000000000000000111111111000000000000000,
    64'b0000000000000000111111111000000000000000111111110000000000000000,
    64'b0000000000000000011111111000000000000000011111110000000000000000,
    64'b0000000000000000011111110000000000000000011111110000000000000000,
    64'b0000000000000000001111110000000000000000011111110000000000000000,
    64'b0000000000000000001111100000000000000000011111100000000000000000,
    64'b0000000000000000001111100000000000000000001111000000000000000000,
    64'b0000000000000000000011000000000000000000001111000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000
};

logic [31:0] i1_bitmap [0:63] = {
    64'b00000000000000000000000000000000,
    64'b00000000000000000000000000000000,
    64'b00000000000000000000000000000000,
    64'b00000000000000000000000000000000,
    64'b00000000000000000000000000000000,
    64'b00000000011111111111110000000000,
    64'b00000001111111111111111000000000,
    64'b00000011111111111111111110000000,
    64'b00000111111100000000111111100000,
    64'b00001111110000000000011111100000,
    64'b00001111100000000000001111110000,
    64'b00001110000000000000000111110000,
    64'b00001110000000000000000111110000,
    64'b00001110000000000000000111110000,
    64'b00001110000000000000000111110000,
    64'b00011110000000000000000111110000,
    64'b00011110000000000000000111110000,
    64'b00011110000000000000000111110000,
    64'b00011110000000000000000111110000,
    64'b00011110000000000000000111110000,
    64'b00011110000000000000000111110000,
    64'b00011110000000000000000111110000,
    64'b00011110000000000000000111110000,
    64'b00011110000000000000000111110000,
    64'b00011110000000000000000111110000,
    64'b00011110000000000000000111110000,
    64'b00011110000000000000000111110000,
    64'b00011110000000000000000111110000,
    64'b00011110000000000000000111110000,
    64'b00011110000000000000000111110000,
    64'b00011110000000000000000111110000,
    64'b00011110000000000000000111110000,
    64'b00011110000000000000000111110000,
    64'b00011110000000000000000111110000,
    64'b00011110000000000000000111110000,
    64'b00011110000000000000000111110000,
    64'b00011110000000000000000111110000,
    64'b00011110000000000000000111110000,
    64'b00011110000000000000000111110000,
    64'b00011110000000000000000111110000,
    64'b00011110000000000000000111110000,
    64'b00011110000000000000000111110000,
    64'b00011110000000000000000111110000,
    64'b00011110000000000000000111110000,
    64'b00011110000000000000000111110000,
    64'b00011110000000000000000111110000,
    64'b00011110000000000000000111110000,
    64'b00011110000000000000000111110000,
    64'b00011110000000000000000111110000,
    64'b00011110000000000000000111110000,
    64'b00011110000000000000000111110000,
    64'b00011110000000000000000111110000,
    64'b00011110000000000000000111110000,
    64'b00011110000000000000000111110000,
    64'b00011110000000000000000111110000,
    64'b00001111100000000000001111110000,
    64'b00000111111111111111111111000000,
    64'b00000011111111111111111110000000,
    64'b00000000011111111111110000000000,
    64'b00000000000011111000000000000000,
    64'b00000000000000000000000000000000,
    64'b00000000000000000000000000000000,
    64'b00000000000000000000000000000000,
    64'b00000000000000000000000000000000
};

logic [31:0] i2_bitmap [0:63] = {
    64'b00000000000000000000000000000000,
    64'b00000000000000000000000000000000,
    64'b00000000000000000000000000000000,
    64'b00000000000000000000000000000000,
    64'b00000000000000000000000000000000,
    64'b00000000000000000000000000000000,
    64'b00000000000000000000000000000000,
    64'b00000000000000000000000000000000,
    64'b00000000111111111111110000000000,
    64'b00000001111111111111111000000000,
    64'b00000001111111111111111000000000,
    64'b00000001111111111111111000000000,
    64'b00000001111111111111111000000000,
    64'b00000001111111111111111000000000,
    64'b00000001111111111111111000000000,
    64'b00000001111111111111111000000000,
    64'b00000001111111111111111000000000,
    64'b00000001111111111111111000000000,
    64'b00000001111111111111111000000000,
    64'b00000001111111111111111000000000,
    64'b00000001111111111111111000000000,
    64'b00000001111111111111111000000000,
    64'b00000001111111111111111000000000,
    64'b00000001111111111111111000000000,
    64'b00000001111111111111111000000000,
    64'b00000001111111111111111000000000,
    64'b00000001111111111111111000000000,
    64'b00000001111111111111111000000000,
    64'b00000001111111111111111000000000,
    64'b00000001111111111111111000000000,
    64'b00000001111111111111111000000000,
    64'b00000001111111111111111000000000,
    64'b00000001111111111111111000000000,
    64'b00000001111111111111111000000000,
    64'b00000001111111111111111000000000,
    64'b00000001111111111111111000000000,
    64'b00000001111111111111111000000000,
    64'b00000001111111111111111000000000,
    64'b00000001111111111111111000000000,
    64'b00000001111111111111111000000000,
    64'b00000001111111111111111000000000,
    64'b00000001111111111111111000000000,
    64'b00000001111111111111111000000000,
    64'b00000001111111111111111000000000,
    64'b00000001111111111111111000000000,
    64'b00000001111111111111111000000000,
    64'b00000001111111111111111000000000,
    64'b00000001111111111111111000000000,
    64'b00000001111111111111111000000000,
    64'b00000001111111111111111000000000,
    64'b00000001111111111111111000000000,
    64'b00000001111111111111111000000000,
    64'b00000001111111111111111000000000,
    64'b00000001111111111111111000000000,
    64'b00000001111111111111111000000000,
    64'b00000000111111111111110000000000,
    64'b00000000000000000000000000000000,
    64'b00000000000000000000000000000000,
    64'b00000000000000000000000000000000,
    64'b00000000000000000000000000000000,
    64'b00000000000000000000000000000000,
    64'b00000000000000000000000000000000,
    64'b00000000000000000000000000000000,
    64'b00000000000000000000000000000000
};

logic [31:0] i3_bitmap [0:63] = {
    64'b00000000000000000000000000000000,
    64'b00000000000000000000000000000000,
    64'b00000000000000000000000000000000,
    64'b00000000000000000000000000000000,
    64'b00000000000000000000000000000000,
    64'b00000000000000000000000000000000,
    64'b00000000000000000000000000000000,
    64'b00000000000000000000000000000000,
    64'b00000000000000000000000000000000,
    64'b00000000000000000000000000000000,
    64'b00000000000000000000000000000000,
    64'b00000000000000000000000000000000,
    64'b00000000000000000000000000000000,
    64'b00000000000111111110000000000000,
    64'b00000000001111111111000000000000,
    64'b00000000001111111111000000000000,
    64'b00000000001111111111000000000000,
    64'b00000000001111111111000000000000,
    64'b00000000001111111111000000000000,
    64'b00000000001111111111000000000000,
    64'b00000000001111111111000000000000,
    64'b00000000001111111111000000000000,
    64'b00000000001111111111000000000000,
    64'b00000000001111111111000000000000,
    64'b00000000001111111111000000000000,
    64'b00000000001111111111000000000000,
    64'b00000000001111111111000000000000,
    64'b00000000001111111111000000000000,
    64'b00000000001111111111000000000000,
    64'b00000000001111111111000000000000,
    64'b00000000001111111111000000000000,
    64'b00000000001111111111000000000000,
    64'b00000000001111111111000000000000,
    64'b00000000001111111111000000000000,
    64'b00000000001111111111000000000000,
    64'b00000000001111111111000000000000,
    64'b00000000001111111111000000000000,
    64'b00000000001111111111000000000000,
    64'b00000000001111111111000000000000,
    64'b00000000001111111111000000000000,
    64'b00000000001111111111000000000000,
    64'b00000000001111111111000000000000,
    64'b00000000001111111111000000000000,
    64'b00000000001111111111000000000000,
    64'b00000000001111111111000000000000,
    64'b00000000001111111111000000000000,
    64'b00000000001111111111000000000000,
    64'b00000000001111111111000000000000,
    64'b00000000001111111111000000000000,
    64'b00000000001111111111000000000000,
    64'b00000000000111111110000000000000,
    64'b00000000000000000000000000000000,
    64'b00000000000000000000000000000000,
    64'b00000000000000000000000000000000,
    64'b00000000000000000000000000000000,
    64'b00000000000000000000000000000000,
    64'b00000000000000000000000000000000,
    64'b00000000000000000000000000000000,
    64'b00000000000000000000000000000000,
    64'b00000000000000000000000000000000,
    64'b00000000000000000000000000000000,
    64'b00000000000000000000000000000000,
    64'b00000000000000000000000000000000,
    64'b00000000000000000000000000000000
};

    logic [31:0] ex1_bitmap [0:63] = {
    64'b00000000000000000000000000000000,
    64'b00000000000000000000000000000000,
    64'b00000000000000000000000000000000,
    64'b00000000000000000000000000000000,
    64'b00000000000000000000000000000000,
    64'b00000000000111111111111100000000,
    64'b00000000011111111111111110000000,
    64'b00000000111111111111111111000000,
    64'b00000011111000000000001111111000,
    64'b00000011110000000000000111111000,
    64'b00001111100000000000000011111100,
    64'b00001111000000000000000001111100,
    64'b00001111000000000000000001111100,
    64'b00001111000000000000000001111100,
    64'b00001111000000000000000001111100,
    64'b00001111000000000000000001111100,
    64'b00001111000000000000000001111100,
    64'b00001111000000000000000001111100,
    64'b00001111000000000000000001111100,
    64'b00001111000000000000000001111100,
    64'b00001111000000000000000001111100,
    64'b00001111000000000000000001111100,
    64'b00001111000000000000000001111100,
    64'b00001111000000000000000001111100,
    64'b00001111000000000000000001111100,
    64'b00001111000000000000000001111100,
    64'b00001111000000000000000001111100,
    64'b00001111000000000000000001111100,
    64'b00001111000000000000000001111100,
    64'b00001111000000000000000001111100,
    64'b00001111000000000000000001111100,
    64'b00001111000000000000000001111100,
    64'b00001111000000000000000001111100,
    64'b00001111000000000000000001111100,
    64'b00001111000000000000000001111100,
    64'b00001111000000000000000001111100,
    64'b00001111000000000000000001111100,
    64'b00001111000000000000000001111100,
    64'b00001111000000000000000001111100,
    64'b00001111000000000000000001111100,
    64'b00001111000000000000000001111100,
    64'b00001111000000000000000001111100,
    64'b00001111000000000000000001111100,
    64'b00001111000000000000000001111100,
    64'b00001111000000000000000001111100,
    64'b00001111000000000000000001111100,
    64'b00001111000000000000000001111100,
    64'b00001111000000000000000001111100,
    64'b00001111000000000000000001111100,
    64'b00001111000000000000000001111100,
    64'b00001111000000000000000001111100,
    64'b00001111000000000000000001111100,
    64'b00001111000000000000000001111100,
    64'b00001111000000000000000001111100,
    64'b00001111100000000000000011111100,
    64'b00000011110000000000000111111000,
    64'b00000001111111111111111111000000,
    64'b00000001111111111111111110000000,
    64'b00000000011111111111111100000000,
    64'b00000000000111111111110000000000,
    64'b00000000000000000000000000000000,
    64'b00000000000000000000000000000000,
    64'b00000000000000000000000000000000,
    64'b00000000000000000000000000000000
};

    logic [31:0] ex2_bitmap [0:63] = {
    64'b00000000000000000000000000000000,
    64'b00000000000000000000000000000000,
    64'b00000000000000000000000000000000,
    64'b00000000000000000000000000000000,
    64'b00000000000000000000000000000000,
    64'b00000000000000000000000000000000,
    64'b00000000000000000000000000000000,
    64'b00000000000000000000000000000000,
    64'b00000000000111111111110000000000,
    64'b00000000001111111111111000000000,
    64'b00000000011111111111111100000000,
    64'b00000000111111111111111110000000,
    64'b00000000111111111111111110000000,
    64'b00000000111111111111111110000000,
    64'b00000000111111111111111110000000,
    64'b00000000111111111111111110000000,
    64'b00000000111111111111111110000000,
    64'b00000000111111111111111110000000,
    64'b00000000111111111111111110000000,
    64'b00000000111111111111111110000000,
    64'b00000000111111111111111110000000,
    64'b00000000111111111111111110000000,
    64'b00000000111111111111111110000000,
    64'b00000000111111111111111110000000,
    64'b00000000111111111111111110000000,
    64'b00000000111111111111111110000000,
    64'b00000000111111111111111110000000,
    64'b00000000111111111111111110000000,
    64'b00000000111111111111111110000000,
    64'b00000000111111111111111110000000,
    64'b00000000111111111111111110000000,
    64'b00000000111111111111111110000000,
    64'b00000000111111111111111110000000,
    64'b00000000111111111111111110000000,
    64'b00000000111111111111111110000000,
    64'b00000000111111111111111110000000,
    64'b00000000111111111111111110000000,
    64'b00000000111111111111111110000000,
    64'b00000000111111111111111110000000,
    64'b00000000111111111111111110000000,
    64'b00000000111111111111111110000000,
    64'b00000000111111111111111110000000,
    64'b00000000111111111111111110000000,
    64'b00000000111111111111111110000000,
    64'b00000000111111111111111110000000,
    64'b00000000111111111111111110000000,
    64'b00000000111111111111111110000000,
    64'b00000000111111111111111110000000,
    64'b00000000111111111111111110000000,
    64'b00000000111111111111111110000000,
    64'b00000000111111111111111110000000,
    64'b00000000111111111111111110000000,
    64'b00000000111111111111111110000000,
    64'b00000000111111111111111110000000,
    64'b00000000011111111111111100000000,
    64'b00000000001111111111111000000000,
    64'b00000000000000000000000000000000,
    64'b00000000000000000000000000000000,
    64'b00000000000000000000000000000000,
    64'b00000000000000000000000000000000,
    64'b00000000000000000000000000000000,
    64'b00000000000000000000000000000000,
    64'b00000000000000000000000000000000,
    64'b00000000000000000000000000000000
};

    logic [31:0] ex3_bitmap [0:63] = {
    64'b00000000000000000000000000000000,
    64'b00000000000000000000000000000000,
    64'b00000000000000000000000000000000,
    64'b00000000000000000000000000000000,
    64'b00000000000000000000000000000000,
    64'b00000000000000000000000000000000,
    64'b00000000000000000000000000000000,
    64'b00000000000000000000000000000000,
    64'b00000000000000000000000000000000,
    64'b00000000000000000000000000000000,
    64'b00000000000000000000000000000000,
    64'b00000000000000000000000000000000,
    64'b00000000000000000000000000000000,
    64'b00000000000000111110000000000000,
    64'b00000000000001111111000000000000,
    64'b00000000000011111111100000000000,
    64'b00000000000011111111100000000000,
    64'b00000000000011111111100000000000,
    64'b00000000000011111111100000000000,
    64'b00000000000011111111100000000000,
    64'b00000000000011111111100000000000,
    64'b00000000000011111111100000000000,
    64'b00000000000011111111100000000000,
    64'b00000000000011111111100000000000,
    64'b00000000000011111111100000000000,
    64'b00000000000011111111100000000000,
    64'b00000000000011111111100000000000,
    64'b00000000000011111111100000000000,
    64'b00000000000011111111100000000000,
    64'b00000000000011111111100000000000,
    64'b00000000000011111111100000000000,
    64'b00000000000011111111100000000000,
    64'b00000000000011111111100000000000,
    64'b00000000000011111111100000000000,
    64'b00000000000011111111100000000000,
    64'b00000000000011111111100000000000,
    64'b00000000000011111111100000000000,
    64'b00000000000011111111100000000000,
    64'b00000000000011111111100000000000,
    64'b00000000000011111111100000000000,
    64'b00000000000001111111000000000000,
    64'b00000000000000111110000000000000,
    64'b00000000000000000000000000000000,
    64'b00000000000000000000000000000000,
    64'b00000000000000000000000000000000,
    64'b00000000000000000000000000000000,
    64'b00000000000000000000000000000000,
    64'b00000000000001111111000000000000,
    64'b00000000000011111111100000000000,
    64'b00000000000011111111100000000000,
    64'b00000000000011111111100000000000,
    64'b00000000000001111111000000000000,
    64'b00000000000000000000000000000000,
    64'b00000000000000000000000000000000,
    64'b00000000000000000000000000000000,
    64'b00000000000000000000000000000000,
    64'b00000000000000000000000000000000,
    64'b00000000000000000000000000000000,
    64'b00000000000000000000000000000000,
    64'b00000000000000000000000000000000,
    64'b00000000000000000000000000000000,
    64'b00000000000000000000000000000000,
    64'b00000000000000000000000000000000,
    64'b00000000000000000000000000000000
};

    logic [63:0] n1_bitmap [0:63] = {
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000011111111110000000000000000000000000000111111100000000000,
    64'b0000000111111111111000000000000000000000000001111111111100000000,
    64'b0000001111111111111100000000000000000000000011111111111110000000,
    64'b0000111111000000111111100000000000000000001111110000001111100000,
    64'b0000111100000000001111110000000000000000011111000000000011100000,
    64'b0000111100000000000111110000000000000000011110000000000011110000,
    64'b0000111000000000000011111000000000000000011110000000000001110000,
    64'b0001110000000000000001111110000000000000011110000000000001110000,
    64'b0001110000000000000000111111000000000000011100000000000001110000,
    64'b0001110000000000000000001111100000000000011100000000000001111000,
    64'b0001110000000000000000001111100000000000011100000000000001111000,
    64'b0001110000000000000000000111110000000000011100000000000001111000,
    64'b0001110000000000000000000011111100000000011100000000000001111000,
    64'b0001110000000000000000000001111110000000011100000000000001111000,
    64'b0001110000000000000000000000111111000000011100000000000001111000,
    64'b0001110000000000000000000000011111100000011100000000000001111000,
    64'b0001110000000000000000000000001111100000011100000000000001111000,
    64'b0001110000000000000000000000000111111000011100000000000001110000,
    64'b0001110000000000000000000000000011111100011100000000000001110000,
    64'b0001110000000000000000000000000000111111011100000000000001111000,
    64'b0001110000000000000000000000000000011111011100000000000001111000,
    64'b0001110000000000000000000000000000001111111100000000000001111000,
    64'b0001110000000000000000000000000000000111111100000000000001111000,
    64'b0001110000000000000000000000000000000011111100000000000001111000,
    64'b0001110000000000000000000000000000000001111100000000000001111000,
    64'b0001110000000000000000000000000000000000111100000000000001111000,
    64'b0001110000000000000100000000000000000000111100000000000001111000,
    64'b0001110000000000000110000000000000000000001100000000000001111000,
    64'b0001110000000000000111000000000000000000000100000000000001111000,
    64'b0001110000000000000111110000000000000000000000000000000001111000,
    64'b0001110000000000000111110000000000000000000000000000000001111000,
    64'b0001110000000000000111111000000000000000000000000000000001111000,
    64'b0001110000000000000111111100000000000000000000000000000001111000,
    64'b0001110000000000000111111110000000000000000000000000000001111000,
    64'b0001110000000000000111011111100000000000000000000000000001111000,
    64'b0001110000000000000111001111110000000000000000000000000001111000,
    64'b0001110000000000000111000011111000000000000000000000000001111000,
    64'b0001110000000000000111000001111110000000000000000000000001111000,
    64'b0001110000000000000111000000111111000000000000000000000001111000,
    64'b0001110000000000000111000000011111100000000000000000000001111000,
    64'b0001110000000000000111000000011111100000000000000000000001111000,
    64'b0001110000000000000111000000000111110000000000000000000001111000,
    64'b0001110000000000000111000000000011111000000000000000000001111000,
    64'b0001110000000000000111000000000001111100000000000000000001111000,
    64'b0001110000000000000111000000000000111111000000000000000001111000,
    64'b0001110000000000000111000000000000011111000000000000000001111000,
    64'b0001110000000000000111000000000000001111100000000000000001111000,
    64'b0001110000000000000111000000000000000111110000000000000001111000,
    64'b0001111000000000000111000000000000000011111100000000000001110000,
    64'b0001111000000000000111000000000000000001111110000000000011110000,
    64'b0001111100000000001111000000000000000000111110000000000011100000,
    64'b0000111111111111111100000000000000000000001111111111111111000000,
    64'b0000011111111111111000000000000000000000000111111111111100000000,
    64'b0000001111111111111000000000000000000000000011111111111000000000,
    64'b0000000011111111100000000000000000000000000001111111100000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000
};

    logic [63:0] n2_bitmap [0:63] = {
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000111111000000000000000000000000000000001111110000000000,
    64'b0000000011111111110000000000000000000000000000111111111100000000,
    64'b0000000011111111111000000000000000000000000001111111111100000000,
    64'b0000000111111111111100000000000000000000000001111111111110000000,
    64'b0000001111111111111110000000000000000000000001111111111110000000,
    64'b0000001111111111111111000000000000000000000011111111111110000000,
    64'b0000001111111111111111110000000000000000000011111111111110000000,
    64'b0000001111111111111111110000000000000000000011111111111110000000,
    64'b0000001111111111111111111000000000000000000011111111111110000000,
    64'b0000001111111111111111111100000000000000000011111111111110000000,
    64'b0000001111111111111111111110000000000000000011111111111110000000,
    64'b0000001111111111111111111111000000000000000011111111111110000000,
    64'b0000001111111111111111111111100000000000000011111111111110000000,
    64'b0000001111111111111111111111110000000000000011111111111110000000,
    64'b0000001111111111111111111111111000000000000011111111111110000000,
    64'b0000001111111111111111111111111100000000000011111111111110000000,
    64'b0000001111111111111111111111111111000000000011111111111110000000,
    64'b0000001111111111111111111111111111100000000011111111111110000000,
    64'b0000001111111111111111111111111111110000000011111111111110000000,
    64'b0000001111111111111111111111111111111000000011111111111110000000,
    64'b0000001111111111111111111111111111111100000011111111111110000000,
    64'b0000001111111111111111111111111111111110000011111111111110000000,
    64'b0000001111111111111111111111111111111111000011111111111110000000,
    64'b0000001111111111111011111111111111111111000011111111111110000000,
    64'b0000001111111111111001111111111111111111110011111111111110000000,
    64'b0000001111111111111000111111111111111111111011111111111110000000,
    64'b0000001111111111111000001111111111111111111111111111111110000000,
    64'b0000001111111111111000001111111111111111111111111111111110000000,
    64'b0000001111111111111000000111111111111111111111111111111110000000,
    64'b0000001111111111111000000011111111111111111111111111111110000000,
    64'b0000001111111111111000000001111111111111111111111111111110000000,
    64'b0000001111111111111000000000011111111111111111111111111110000000,
    64'b0000001111111111111000000000001111111111111111111111111110000000,
    64'b0000001111111111111000000000000111111111111111111111111110000000,
    64'b0000001111111111111000000000000001111111111111111111111110000000,
    64'b0000001111111111111000000000000000111111111111111111111110000000,
    64'b0000001111111111111000000000000000011111111111111111111110000000,
    64'b0000001111111111111000000000000000011111111111111111111110000000,
    64'b0000001111111111111000000000000000001111111111111111111110000000,
    64'b0000001111111111111000000000000000000111111111111111111110000000,
    64'b0000001111111111111000000000000000000011111111111111111110000000,
    64'b0000001111111111111000000000000000000000111111111111111110000000,
    64'b0000001111111111111000000000000000000000111111111111111110000000,
    64'b0000001111111111111000000000000000000000011111111111111110000000,
    64'b0000001111111111111000000000000000000000001111111111111110000000,
    64'b0000001111111111111000000000000000000000000011111111111110000000,
    64'b0000000111111111111000000000000000000000000001111111111110000000,
    64'b0000000011111111110000000000000000000000000001111111111110000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000
};

    logic [63:0] n3_bitmap [0:63] = {
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000111111100000000000000000000000000000001111110000000000,
    64'b0000000000111111100000000000000000000000000000001111110000000000,
    64'b0000000000111111110000000000000000000000000000001111110000000000,
    64'b0000000000111111111000000000000000000000000000001111110000000000,
    64'b0000000000111111111100000000000000000000000000001111110000000000,
    64'b0000000000111111111110000000000000000000000000001111110000000000,
    64'b0000000000111111111111000000000000000000000000001111110000000000,
    64'b0000000000111111111111100000000000000000000000001111110000000000,
    64'b0000000000111111111111111000000000000000000000001111110000000000,
    64'b0000000000111111111111111000000000000000000000001111110000000000,
    64'b0000000000111111111111111100000000000000000000001111110000000000,
    64'b0000000000111111111111111110000000000000000000001111110000000000,
    64'b0000000000111111001111111111100000000000000000001111110000000000,
    64'b0000000000111111000111111111100000000000000000001111110000000000,
    64'b0000000000111111000011111111111000000000000000001111110000000000,
    64'b0000000000111111000000111111111100000000000000001111110000000000,
    64'b0000000000111111000000111111111110000000000000001111110000000000,
    64'b0000000000111111000000011111111111000000000000001111110000000000,
    64'b0000000000111111000000001111111111100000000000001111110000000000,
    64'b0000000000111111000000000111111111100000000000001111110000000000,
    64'b0000000000111111000000000011111111111000000000001111110000000000,
    64'b0000000000111111000000000000111111111100000000001111110000000000,
    64'b0000000000111111000000000000011111111110000000001111110000000000,
    64'b0000000000111111000000000000011111111111000000001111110000000000,
    64'b0000000000111111000000000000001111111111100000001111110000000000,
    64'b0000000000111111000000000000000011111111110000001111110000000000,
    64'b0000000000111111000000000000000001111111110000001111110000000000,
    64'b0000000000111111000000000000000000111111111100001111110000000000,
    64'b0000000000111111000000000000000000011111111111001111110000000000,
    64'b0000000000111111000000000000000000000111111111101111110000000000,
    64'b0000000000111111000000000000000000000011111111111111110000000000,
    64'b0000000000111111000000000000000000000001111111111111110000000000,
    64'b0000000000111111000000000000000000000000111111111111110000000000,
    64'b0000000000111111000000000000000000000000011111111111110000000000,
    64'b0000000000111111000000000000000000000000001111111111110000000000,
    64'b0000000000111111000000000000000000000000000111111111110000000000,
    64'b0000000000111111000000000000000000000000000011111111110000000000,
    64'b0000000000111111000000000000000000000000000001111111110000000000,
    64'b0000000000111111000000000000000000000000000000111111110000000000,
    64'b0000000000111111000000000000000000000000000000011111110000000000,
    64'b0000000000111111000000000000000000000000000000001111110000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000
};

logic [63:0] Lout_bitmap [0:63] = {
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000011111111111110000000000000000000000000000000000000000,
    64'b0000000000111111111111111000000000000000000000000000000000000000,
    64'b0000000001111111111111111100000000000000000000000000000000000000,
    64'b0000000001111100000000111110000000000000000000000000000000000000,
    64'b0000000001111000000000111111000000000000000000000000000000000000,
    64'b0000000011110000000000011111000000000000000000000000000000000000,
    64'b0000000011110000000000001111000000000000000000000000000000000000,
    64'b0000000011110001111110000111000000000000000000000000000000000000,
    64'b0000000011100011111111000111000000000000000000000000000000000000,
    64'b0000000011100011111111000111000000000000000000000000000000000000,
    64'b0000000011100011111111000111000000000000000000000000000000000000,
    64'b0000000011100011100111000111000000000000000000000000000000000000,
    64'b0000000011100011100111000111000000000000000000000000000000000000,
    64'b0000000011100011100111000111000000000000000000000000000000000000,
    64'b0000000011100011100111000111000000000000000000000000000000000000,
    64'b0000000011100011100111000111000000000000000000000000000000000000,
    64'b0000000011100011100111000111000000000000000000000000000000000000,
    64'b0000000011100011100111000111000000000000000000000000000000000000,
    64'b0000000011100011100111000111000000000000000000000000000000000000,
    64'b0000000011100011100111000111000000000000000000000000000000000000,
    64'b0000000011100011100111000111000000000000000000000000000000000000,
    64'b0000000011100011100111000111000000000000000000000000000000000000,
    64'b0000000011100011100111000111000000000000000000000000000000000000,
    64'b0000000011100011100111000111000000000000000000000000000000000000,
    64'b0000000011100011100111000111000000000000000000000000000000000000,
    64'b0000000011100011100111000111000000000000000000000000000000000000,
    64'b0000000011100011100111000111000000000000000000000000000000000000,
    64'b0000000011100011100111000111000000000000000000000000000000000000,
    64'b0000000011100011100111000111000000000000000000000000000000000000,
    64'b0000000011100011100111000111000000000000000000000000000000000000,
    64'b0000000011100011100111000111000000000000000000000000000000000000,
    64'b0000000011100011100111000111000000000000000000000000000000000000,
    64'b0000000011100011100111000111000000000000000000000000000000000000,
    64'b0000000011100011100111000111000000000000000000000000000000000000,
    64'b0000000011100011100111000111000000000000000000000000000000000000,
    64'b0000000011100011110111000111110000000000000000000000000000000000,
    64'b0000000011100011110111000111111100000000000000000000000000000000,
    64'b0000000011100011110111111111111111111111111111111111111110000000,
    64'b0000000011100001110111111111111111111111111111111111111111100000,
    64'b0000000011100001111111111111111111111111111111111111111111110000,
    64'b0000000011110001111111111111111111111111111110000000001111111000,
    64'b0000000011110001111111111111111111111110000000000000000011111000,
    64'b0000000011110000111111111100000000000000000000000000000001111000,
    64'b0000000001110000111111111111111111111111111111111111110000111000,
    64'b0000000001110000011111111111111111111111111111111111111000111000,
    64'b0000000001110000011111111111111111111111111111111111111000111000,
    64'b0000000001111000000111111111111111111111111111111111111000111000,
    64'b0000000001111100000001111111111111111111111111111111111000111000,
    64'b0000000001111110000000001111111111111111111111111111110000111000,
    64'b0000000000111111000000000000000000000000000000000000000000111000,
    64'b0000000000011111100000000000000000000000000000000000000000111000,
    64'b0000000000001111110000000000000000000000000000000000000001111000,
    64'b0000000000000111111111000000000000000000000000000000000001111000,
    64'b0000000000000011111111111111111111111111111111111111111111111000,
    64'b0000000000000001111111111111111111111111111111111111111111110000,
    64'b0000000000000000000111111111111111111111111111111111111111110000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000
};



logic [63:0] Lmid_bitmap [0:63] = {
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000011111111000000000000000000000000000000000000000000,
    64'b0000000000000111111111000000000000000000000000000000000000000000,
    64'b0000000000001111111111100000000000000000000000000000000000000000,
    64'b0000000000001111111111110000000000000000000000000000000000000000,
    64'b0000000000001110000001111000000000000000000000000000000000000000,
    64'b0000000000011100000000111000000000000000000000000000000000000000,
    64'b0000000000011100000000111000000000000000000000000000000000000000,
    64'b0000000000011100000000111000000000000000000000000000000000000000,
    64'b0000000000011100000000111000000000000000000000000000000000000000,
    64'b0000000000011100000000111000000000000000000000000000000000000000,
    64'b0000000000011100000000111000000000000000000000000000000000000000,
    64'b0000000000011100000000111000000000000000000000000000000000000000,
    64'b0000000000011100000000111000000000000000000000000000000000000000,
    64'b0000000000011100000000111000000000000000000000000000000000000000,
    64'b0000000000011100000000111000000000000000000000000000000000000000,
    64'b0000000000011100000000111000000000000000000000000000000000000000,
    64'b0000000000011100000000111000000000000000000000000000000000000000,
    64'b0000000000011100000000111000000000000000000000000000000000000000,
    64'b0000000000011100000000111000000000000000000000000000000000000000,
    64'b0000000000011100000000111000000000000000000000000000000000000000,
    64'b0000000000011100000000111000000000000000000000000000000000000000,
    64'b0000000000011100000000111000000000000000000000000000000000000000,
    64'b0000000000011100000000111000000000000000000000000000000000000000,
    64'b0000000000011100000000111000000000000000000000000000000000000000,
    64'b0000000000011100000000111000000000000000000000000000000000000000,
    64'b0000000000011100000000111000000000000000000000000000000000000000,
    64'b0000000000011100000000111000000000000000000000000000000000000000,
    64'b0000000000011100000000111000000000000000000000000000000000000000,
    64'b0000000000011100000000111000000000000000000000000000000000000000,
    64'b0000000000011100000000111000000000000000000000000000000000000000,
    64'b0000000000011100000000111000000000000000000000000000000000000000,
    64'b0000000000011100000000111000000000000000000000000000000000000000,
    64'b0000000000011100000000111000000000000000000000000000000000000000,
    64'b0000000000011100000000111000000000000000000000000000000000000000,
    64'b0000000000011100000000111000000000000000000000000000000000000000,
    64'b0000000000011110000000111100000000000000000000000000000000000000,
    64'b0000000000011110000000111110000000000000000000000000000000000000,
    64'b0000000000001110000000111111111111111111111111111111110000000000,
    64'b0000000000001110000000011111111111111111111111111111111100000000,
    64'b0000000000001111000000000011111111111111111111111111111110000000,
    64'b0000000000001111000000000000000000000000000000000000001111000000,
    64'b0000000000001111100000000000000000000000000000000000000111000000,
    64'b0000000000001111100000000000000000000000000000000000000111000000,
    64'b0000000000000111111000000000000000000000000000000000000111000000,
    64'b0000000000000011111110000000000000000000000000000000000111000000,
    64'b0000000000000001111111110000000000000000000000000000001111000000,
    64'b0000000000000000111111111111111111111111111111111111111111000000,
    64'b0000000000000000011111111111111111111111111111111111111111000000,
    64'b0000000000000000001111111111111111111111111111111111111110000000,
    64'b0000000000000000000000111111111111111111111111111111111110000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000
};


logic [63:0] Lin_bitmap [0:63] = {
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000001111110000000000000000000000000000000000000000000,
    64'b0000000000000011111111000000000000000000000000000000000000000000,
    64'b0000000000000011111111000000000000000000000000000000000000000000,
    64'b0000000000000011111111000000000000000000000000000000000000000000,
    64'b0000000000000011111111000000000000000000000000000000000000000000,
    64'b0000000000000011111111000000000000000000000000000000000000000000,
    64'b0000000000000011111111000000000000000000000000000000000000000000,
    64'b0000000000000011111111000000000000000000000000000000000000000000,
    64'b0000000000000011111111000000000000000000000000000000000000000000,
    64'b0000000000000011111111000000000000000000000000000000000000000000,
    64'b0000000000000011111111000000000000000000000000000000000000000000,
    64'b0000000000000011111111000000000000000000000000000000000000000000,
    64'b0000000000000011111111000000000000000000000000000000000000000000,
    64'b0000000000000011111111000000000000000000000000000000000000000000,
    64'b0000000000000011111111000000000000000000000000000000000000000000,
    64'b0000000000000011111111000000000000000000000000000000000000000000,
    64'b0000000000000011111111000000000000000000000000000000000000000000,
    64'b0000000000000011111111000000000000000000000000000000000000000000,
    64'b0000000000000011111111000000000000000000000000000000000000000000,
    64'b0000000000000011111111000000000000000000000000000000000000000000,
    64'b0000000000000011111111000000000000000000000000000000000000000000,
    64'b0000000000000011111111000000000000000000000000000000000000000000,
    64'b0000000000000011111111000000000000000000000000000000000000000000,
    64'b0000000000000011111111000000000000000000000000000000000000000000,
    64'b0000000000000011111111000000000000000000000000000000000000000000,
    64'b0000000000000011111111000000000000000000000000000000000000000000,
    64'b0000000000000011111111000000000000000000000000000000000000000000,
    64'b0000000000000011111111000000000000000000000000000000000000000000,
    64'b0000000000000011111111000000000000000000000000000000000000000000,
    64'b0000000000000011111111000000000000000000000000000000000000000000,
    64'b0000000000000011111111000000000000000000000000000000000000000000,
    64'b0000000000000001111111000000000000000000000000000000000000000000,
    64'b0000000000000001111111000000000000000000000000000000000000000000,
    64'b0000000000000001111111000000000000000000000000000000000000000000,
    64'b0000000000000001111111100000000000000000000000000000000000000000,
    64'b0000000000000000111111111100000000000000000000000000000000000000,
    64'b0000000000000000111111111111111111111111111111111111110000000000,
    64'b0000000000000000011111111111111111111111111111111111111000000000,
    64'b0000000000000000011111111111111111111111111111111111111000000000,
    64'b0000000000000000000111111111111111111111111111111111111000000000,
    64'b0000000000000000000001111111111111111111111111111111111000000000,
    64'b0000000000000000000000001111111111111111111111111111110000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000
};

// 이거 안에 검정 테두리가 없음 나중에 수정해봐 
/***************************/
logic [63:0] Oout_bitmap[0:63] = {
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000111111111111111111111111111111100000000000000000,
    64'b0000000000001111111111111111111111111111111111111111000000000000,
    64'b0000000000111111111111111111111111111111111111111111110000000000,
    64'b0000000011111111111000000000000000000000000011111111111000000000,
    64'b0000000111111110000000000000000000000000000000000111111100000000,
    64'b0000001111111000000000000000000000000000000000000001111110000000,
    64'b0000011111100000000000000000000000000000000000000000111111000000,
    64'b0000011111000000000000000000000000000000000000000000011111000000,
    64'b0000011110000000000000000000000000000000000000000000001111100000,
    64'b0000111100000000000000000000000000000000000000000000000111100000,
    64'b0000111100000000000000000000000000000000000000000000000111100000,
    64'b0001111100000000000000000000000000000000000000000000000011100000,
    64'b0001111000000000000000000000000000000000000000000000000011100000,
    64'b0001111000000000000000000000000000000000000000000000000011100000,
    64'b0001110000000000000000000000000000000000000000000000000011100000,
    64'b0001110000000000000000000000000000000000000000000000000011100000,
    64'b0001110000000000000000000000000000000000000000000000000011100000,
    64'b0001110000000000000000000000000000000000000000000000000011100000,
    64'b0001110000000000000000011111111111111111000000000000000011100000,
    64'b0001110000000000000011111111111111111111110000000000000011100000,
    64'b0001110000000000000111111111111111111111111000000000000011100000,
    64'b0001110000000000000111111100000000000111111000000000000011100000,
    64'b0001110000000000000111100000000000000001111000000000000011100000,
    64'b0001110000000000000111000000000000000000111000000000000011100000,
    64'b0001110000000000000111000000000000000000111000000000000011100000,
    64'b0001110000000000000111000000000000000000111000000000000011100000,
    64'b0001110000000000000111000000000000000000111000000000000011100000,
    64'b0001110000000000000111000000000000000000111000000000000011100000,
    64'b0001110000000000000111000000000000000000111000000000000011100000,
    64'b0001110000000000000111000000000000000000111000000000000011100000,
    64'b0001110000000000000111000000000000000000111000000000000011100000,
    64'b0001110000000000000111000000000000000000111000000000000011100000,
    64'b0001110000000000000111000000000000000000111000000000000011100000,
    64'b0001110000000000000111000000000000000000111000000000000011100000,
    64'b0001110000000000000111100000000000000001111000000000000011100000,
    64'b0001110000000000000111111110000000000111111000000000000011100000,
    64'b0001110000000000000111111111111111111111111000000000000011100000,
    64'b0001110000000000000011111111111111111111110000000000000011100000,
    64'b0001110000000000000000001111111111111111000000000000000011100000,
    64'b0001110000000000000000000000000000000000000000000000000011100000,
    64'b0001110000000000000000000000000000000000000000000000000011100000,
    64'b0001110000000000000000000000000000000000000000000000000011100000,
    64'b0001111000000000000000000000000000000000000000000000000011100000,
    64'b0001111000000000000000000000000000000000000000000000000011100000,
    64'b0001111000000000000000000000000000000000000000000000000011100000,
    64'b0000111100000000000000000000000000000000000000000000000011100000,
    64'b0000111100000000000000000000000000000000000000000000000111100000,
    64'b0000111110000000000000000000000000000000000000000000001111100000,
    64'b0000011111000000000000000000000000000000000000000000011111100000,
    64'b0000011111100000000000000000000000000000000000000000111111000000,
    64'b0000001111111000000000000000000000000000000000000001111110000000,
    64'b0000000111111100000000000000000000000000000000000111111100000000,
    64'b0000000011111111100000000000000000000000000001111111111000000000,
    64'b0000000000111111111111111111111111111111111111111111110000000000,
    64'b0000000000011111111111111111111111111111111111111111000000000000,
    64'b0000000000000011111111111111111111111111111111110000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000
};


logic [63:0] Omid_bitmap [0:63] = {
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000111111111111111111111111100000000000000000000,
    64'b0000000000000001111111111111111111111111111111111000000000000000,
    64'b0000000000000111111111111111111111111111111111111110000000000000,
    64'b0000000000011111111111111111111111111111111111111111000000000000,
    64'b0000000000111111111110000000000000000000000111111111100000000000,
    64'b0000000001111111100000000000000000000000000000011111110000000000,
    64'b0000000011111100000000000000000000000000000000000111111000000000,
    64'b0000000011111000000000000000000000000000000000000001111000000000,
    64'b0000000011110000000000000000000000000000000000000001111100000000,
    64'b0000000111100000000000000000000000000000000000000000111100000000,
    64'b0000000111000000000000000000000000000000000000000000111100000000,
    64'b0000001111000000000001111111111111111111100000000000011100000000,
    64'b0000001110000000000111111111111111111111111100000000011100000000,
    64'b0000001110000000001111111111111111111111111110000000011100000000,
    64'b0000001110000000011111111111111111111111111110000000011100000000,
    64'b0000001110000000011111100000000000000000111111000000011100000000,
    64'b0000001110000000111100000000000000000000001111000000011100000000,
    64'b0000001110000000111000000000000000000000000111000000011100000000,
    64'b0000001110000000111000000000000000000000000111000000011100000000,
    64'b0000001110000000111000000000000000000000000111000000011100000000,
    64'b0000001110000000111000000000000000000000000111000000011100000000,
    64'b0000001110000000111000000000000000000000000111000000011100000000,
    64'b0000001110000000111000000000000000000000000111000000011100000000,
    64'b0000001110000000111000000000000000000000000111000000011100000000,
    64'b0000001110000000111000000000000000000000000111000000011100000000,
    64'b0000001110000000111000000000000000000000000111000000011100000000,
    64'b0000001110000000111000000000000000000000000111000000011100000000,
    64'b0000001110000000111000000000000000000000000111000000011100000000,
    64'b0000001110000000111000000000000000000000000111000000011100000000,
    64'b0000001110000000111000000000000000000000000111000000011100000000,
    64'b0000001110000000111000000000000000000000000111000000011100000000,
    64'b0000001110000000111000000000000000000000000111000000011100000000,
    64'b0000001110000000111000000000000000000000000111000000011100000000,
    64'b0000001110000000111000000000000000000000000111000000011100000000,
    64'b0000001110000000111100000000000000000000001111000000011100000000,
    64'b0000001110000000111111110000000000000000111111000000011100000000,
    64'b0000001110000000011111111111111111111111111111000000011100000000,
    64'b0000001111000000011111111111111111111111111110000000011100000000,
    64'b0000001111000000000111111111111111111111111110000000111100000000,
    64'b0000000111100000000011111111111111111111110000000000111100000000,
    64'b0000000111100000000000000000000000000000000000000001111100000000,
    64'b0000000111110000000000000000000000000000000000000001111100000000,
    64'b0000000011111000000000000000000000000000000000000011111100000000,
    64'b0000000011111100000000000000000000000000000000011111111000000000,
    64'b0000000001111111100000000000000000000000000001111111110000000000,
    64'b0000000000111111111100000000000000000000001111111111100000000000,
    64'b0000000000011111111111111111111111111111111111111111000000000000,
    64'b0000000000000111111111111111111111111111111111111110000000000000,
    64'b0000000000000011111111111111111111111111111111111000000000000000,
    64'b0000000000000000011111111111111111111111111110000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000
};

logic [63:0] Oin_bitmap [0:63] = {
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000001111111111111111111111000000000000000000000,
    64'b0000000000000000011111111111111111111111111111100000000000000000,
    64'b0000000000000011111111111111111111111111111111111000000000000000,
    64'b0000000000000111111111111111111111111111111111111110000000000000,
    64'b0000000000001111111111111111111111111111111111111110000000000000,
    64'b0000000000011111111111111111111111111111111111111111000000000000,
    64'b0000000000111111111111111111111111111111111111111111000000000000,
    64'b0000000000111111111110000000000000000000011111111111100000000000,
    64'b0000000001111111111000000000000000000000000011111111100000000000,
    64'b0000000001111111110000000000000000000000000001111111100000000000,
    64'b0000000001111111100000000000000000000000000001111111100000000000,
    64'b0000000001111111100000000000000000000000000000111111100000000000,
    64'b0000000001111111000000000000000000000000000000111111100000000000,
    64'b0000000001111111100000000000000000000000000000111111100000000000,
    64'b0000000001111111000000000000000000000000000000111111100000000000,
    64'b0000000001111111000000000000000000000000000000111111100000000000,
    64'b0000000001111111000000000000000000000000000000111111100000000000,
    64'b0000000001111111000000000000000000000000000000111111100000000000,
    64'b0000000001111111000000000000000000000000000000111111100000000000,
    64'b0000000001111111000000000000000000000000000000111111100000000000,
    64'b0000000001111111000000000000000000000000000000111111100000000000,
    64'b0000000001111111000000000000000000000000000000111111100000000000,
    64'b0000000001111111000000000000000000000000000000111111100000000000,
    64'b0000000001111111000000000000000000000000000000111111100000000000,
    64'b0000000001111111000000000000000000000000000000111111100000000000,
    64'b0000000001111111000000000000000000000000000000111111100000000000,
    64'b0000000001111111000000000000000000000000000000111111100000000000,
    64'b0000000001111111000000000000000000000000000000111111100000000000,
    64'b0000000001111111000000000000000000000000000000111111100000000000,
    64'b0000000001111111000000000000000000000000000000111111100000000000,
    64'b0000000001111111000000000000000000000000000000111111100000000000,
    64'b0000000001111111000000000000000000000000000000111111100000000000,
    64'b0000000001111111100000000000000000000000000000111111100000000000,
    64'b0000000000111111100000000000000000000000000001111111100000000000,
    64'b0000000000111111111000000000000000000000000001111111000000000000,
    64'b0000000000011111111100000000000000000000001111111111000000000000,
    64'b0000000000011111111111111111111111111111111111111110000000000000,
    64'b0000000000001111111111111111111111111111111111111110000000000000,
    64'b0000000000000111111111111111111111111111111111111100000000000000,
    64'b0000000000000011111111111111111111111111111111000000000000000000,
    64'b0000000000000000011111111111111111111111111110000000000000000000,
    64'b0000000000000000000011111111111111111111110000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000
};

logic [63:0] Sout_bitmap [0:63] = {
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000011111111111111111111000000000000000000000000000,
    64'b0000000000001111111111111111111111111100000000000000000000000000,
    64'b0000000000111111111111111111111111111110000000000000000000000000,
    64'b0000000001111111111100000000000000111110000000000000000000000000,
    64'b0000000011111110000000000000000000011110000000000000000000000000,
    64'b0000000111111000000000000000000000001111000000000000000000000000,
    64'b0000001111110000000000000000000000001111000000000000000000000000,
    64'b0000011111100000000011111111111110001111000000000000000000000000,
    64'b0000011111000000011111111111111110000111000000000000000000000000,
    64'b0000111110000011111111111111111111000111000000000000000000000000,
    64'b0000111100000111111111100000001111000111000000000000000000000000,
    64'b0000111100001111111111111111111111000111000000000000000000000000,
    64'b0001111000001111111111111111111110000111000000000000000000000000,
    64'b0001111000011111111111111111111110001111000000000000000000000000,
    64'b0001111000011111111111100000000000001111000000000000000000000000,
    64'b0001110000011111111100000000000000001111000000000000000000000000,
    64'b0001110000011101111000000000000000011110000000000000000000000000,
    64'b0001110000111101110000000000000000111110000000000000000000000000,
    64'b0001110000111101110000001111111111111111111111100000000000000000,
    64'b0001110000111101110001111111111111111111111111111110000000000000,
    64'b0001110000111001110000111111111111111111111111111111110000000000,
    64'b0001110000111101110000000000000000000000000011111111111000000000,
    64'b0001110000111101110000000000000000000000000000001111111100000000,
    64'b0001110000111111111000000000000000000000000000000001111110000000,
    64'b0001111000011111111110000000000000000000000000000000111111000000,
    64'b0001111000011111111111111111111111111111111100000000011111100000,
    64'b0001111000001111111111111111111111111111111111100000001111110000,
    64'b0000111000001111111111111111111111111111111111111000000111110000,
    64'b0000111100000111111111111111111111111111111111111110000011110000,
    64'b0000111111000000011111111111111111111111111111111111000001110000,
    64'b0000111111100000000000111111111111111111111111111111000001110000,
    64'b0000011111110000000000000000000000000000001111111111100001110000,
    64'b0000000111111000000000000000000000000000000011111111100001110000,
    64'b0000000011111110000000000000000000000000000000111111100001110000,
    64'b0000000001111111111111000000000000000000000000111011100001110000,
    64'b0000000000111111111111111111111111111111100000111011110001110000,
    64'b0000001111111111111111111111111111111111111000111011100001110000,
    64'b0000011111111111111111111111111111111111111000111011100001110000,
    64'b0000111111111111111111111111111111111111000000111011100001110000,
    64'b0000111110000000000000000000000000000000000000111011100001110000,
    64'b0000111100000000000000000000000000000000000000111111100001110000,
    64'b0000111000000000000000000000000000000000000001111111100001110000,
    64'b0000111000000000000000000000000000000000000111111111100001110000,
    64'b0000111000001111111111111111111111111111111111111111000001110000,
    64'b0000111000011111111111111111111111111111111111111111000001110000,
    64'b0000111000011111111111111111111111111111111111111111000001110000,
    64'b0000111000011111111111111111111111111111111111111100000011110000,
    64'b0000111000011111111111111111111111111111111111110000000111110000,
    64'b0000111000001111111111111111111111111111111100000000001111110000,
    64'b0000111000000000000000000000000000000000000000000000011111100000,
    64'b0000111000000000000000000000000000000000000000000000111111000000,
    64'b0000111100000000000000000000000000000000000000000001111110000000,
    64'b0000111110000000000000000000000000000000000000011111111100000000,
    64'b0000111111111111111111111111111111111111111111111111111000000000,
    64'b0000011111111111111111111111111111111111111111111111110000000000,
    64'b0000001111111111111111111111111111111111111111111100000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000
};

logic [63:0] Smid_bitmap [0:63] = {
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000011111111111111000000000000000000000000000000,
    64'b0000000000000001111111111111111111100000000000000000000000000000,
    64'b0000000000000111111111111111111111110000000000000000000000000000,
    64'b0000000000001111111111111111111111110000000000000000000000000000,
    64'b0000000000011111111100000000000001110000000000000000000000000000,
    64'b0000000000111111100000000000000001111000000000000000000000000000,
    64'b0000000001111100000000000000000000111000000000000000000000000000,
    64'b0000000011111000000000000000000000111000000000000000000000000000,
    64'b0000000011110000000000000000000000111000000000000000000000000000,
    64'b0000000111110000000000000000000001111000000000000000000000000000,
    64'b0000000111100000000000000000000001110000000000000000000000000000,
    64'b0000000111100000000000011111111111110000000000000000000000000000,
    64'b0000001111100000000011111111111111110000000000000000000000000000,
    64'b0000001111100000000111111111111111100000000000000000000000000000,
    64'b0000001111000000001111111111111111000000000000000000000000000000,
    64'b0000001111000000001111110000000000000000000000000000000000000000,
    64'b0000001111000000001110000000000000000000000000000000000000000000,
    64'b0000001111000000001111000000000000000000000000000000000000000000,
    64'b0000001111000000001111111111111111111111111100000000000000000000,
    64'b0000001111000000001111111111111111111111111111110000000000000000,
    64'b0000001111000000000111111111111111111111111111111110000000000000,
    64'b0000000111100000000001111111111111111111111111111111000000000000,
    64'b0000000111100000000000000000000000000000000011111111100000000000,
    64'b0000000111110000000000000000000000000000000000011111110000000000,
    64'b0000000111110000000000000000000000000000000000000111111000000000,
    64'b0000000011111000000000000000000000000000000000000001111100000000,
    64'b0000000000111111100000000000000000000000000000000000111110000000,
    64'b0000000000011111111111000000000000000000000000000000111110000000,
    64'b0000000000001111111111111111111111111111110000000000011110000000,
    64'b0000000000000111111111111111111111111111111100000000011110000000,
    64'b0000000000000001111111111111111111111111111111000000011110000000,
    64'b0000000000000000000000111111111111111111111111000000011110000000,
    64'b0000000000000000000000000000000000000000011111000000001110000000,
    64'b0000000000000000000000000000000000000000000111000000011110000000,
    64'b0000000000000000000000000000000000000000000111000000011110000000,
    64'b0000000000000000000000000000000000000000111111000000011110000000,
    64'b0000000001111111111111111111111111111111111111000000011110000000,
    64'b0000000011111111111111111111111111111111111111000000011110000000,
    64'b0000000111111111111111111111111111111111111110000000011110000000,
    64'b0000000111111111111111111111111111111111111000000000011110000000,
    64'b0000000111110000000000000000000000000000000000000000111110000000,
    64'b0000000111100000000000000000000000000000000000000000111110000000,
    64'b0000000111100000000000000000000000000000000000000000111110000000,
    64'b0000000111100000000000000000000000000000000000000011111100000000,
    64'b0000000111100000000000000000000000000000000000001111111000000000,
    64'b0000000111110000000000000000000000000000000011111111110000000000,
    64'b0000000111111111111111111111111111111111111111111111100000000000,
    64'b0000000111111111111111111111111111111111111111111111000000000000,
    64'b0000000011111111111111111111111111111111111111111110000000000000,
    64'b0000000001111111111111111111111111111111111111100000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000
};


logic [63:0] Sin_bitmap [0:63] = {
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000011111111111110000000000000000000000000000000,
    64'b0000000000000000011111111111111110000000000000000000000000000000,
    64'b0000000000000011111111111111111111000000000000000000000000000000,
    64'b0000000000000111111111111111111111000000000000000000000000000000,
    64'b0000000000001111111111111111111111000000000000000000000000000000,
    64'b0000000000001111111111111111111110000000000000000000000000000000,
    64'b0000000000011111111111111111111110000000000000000000000000000000,
    64'b0000000000011111111111100000000000000000000000000000000000000000,
    64'b0000000000011111111100000000000000000000000000000000000000000000,
    64'b0000000000011111111000000000000000000000000000000000000000000000,
    64'b0000000000111111110000000000000000000000000000000000000000000000,
    64'b0000000000111111110000000000000000000000000000000000000000000000,
    64'b0000000000111111110000000000000000000000000000000000000000000000,
    64'b0000000000111111110000000000000000000000000000000000000000000000,
    64'b0000000000111111110000000000000000000000000000000000000000000000,
    64'b0000000000111111110000000000000000000000000000000000000000000000,
    64'b0000000000111111111000000000000000000000000000000000000000000000,
    64'b0000000000011111111110000000000000000000000000000000000000000000,
    64'b0000000000011111111111111111111111111111111100000000000000000000,
    64'b0000000000001111111111111111111111111111111111100000000000000000,
    64'b0000000000001111111111111111111111111111111111111000000000000000,
    64'b0000000000000111111111111111111111111111111111111110000000000000,
    64'b0000000000000000011111111111111111111111111111111111000000000000,
    64'b0000000000000000000000111111111111111111111111111111000000000000,
    64'b0000000000000000000000000000000000000000001111111111100000000000,
    64'b0000000000000000000000000000000000000000000011111111100000000000,
    64'b0000000000000000000000000000000000000000000000111111100000000000,
    64'b0000000000000000000000000000000000000000000000111111100000000000,
    64'b0000000000000000000000000000000000000000000000111111100000000000,
    64'b0000000000000000000000000000000000000000000000111111100000000000,
    64'b0000000000000000000000000000000000000000000000111111100000000000,
    64'b0000000000000000000000000000000000000000000000111111100000000000,
    64'b0000000000000000000000000000000000000000000000111111100000000000,
    64'b0000000000000000000000000000000000000000000000111111100000000000,
    64'b0000000000000000000000000000000000000000000001111111100000000000,
    64'b0000000000000000000000000000000000000000000111111111100000000000,
    64'b0000000000001111111111111111111111111111111111111111000000000000,
    64'b0000000000011111111111111111111111111111111111111111000000000000,
    64'b0000000000011111111111111111111111111111111111111111000000000000,
    64'b0000000000011111111111111111111111111111111111111100000000000000,
    64'b0000000000011111111111111111111111111111111111110000000000000000,
    64'b0000000000001111111111111111111111111111111100000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000
};

logic [63:0] Eout_bitmap [0:63] = {
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000011111111111111111111111000000000000000000000000,
    64'b0000000000001111111111111111111111111111100000000000000000000000,
    64'b0000000000011111111111111111111111111111110000000000000000000000,
    64'b0000000001111111111100000000000000000111111000000000000000000000,
    64'b0000000011111110000000000000000000000011111100000000000000000000,
    64'b0000000111111100000000000000000000000001111100000000000000000000,
    64'b0000001111110000000000000000000000000000111100000000000000000000,
    64'b0000011111100000000011111111111111110000111100000000000000000000,
    64'b0000011111000000111111111111111111110000111110000000000000000000,
    64'b0000111110000001111111111111111111110000111110000000000000000000,
    64'b0001111100000011111111100000000001110000111110000000000000000000,
    64'b0001111100000111111011111111111111110011111110000000000000000000,
    64'b0001111000001111111111111111111111110000111110000000000000000000,
    64'b0001110000011111111111111111111111110000111110000000000000000000,
    64'b0001110000111111111111100000000000000000111110000000000000000000,
    64'b0001110000111111111100000000000000000001111000000000000000000000,
    64'b0001110001111111111000000000000000000011111000000000000000000000,
    64'b0001111000111011111000000000000000000111111000000000000000000000,
    64'b0001110000111011100000001111111111111111110000000000000000000000,
    64'b0001110000111011100001111111111111111111111111111111111111000000,
    64'b0001110000111011100001111111111111111111111111111111111111100000,
    64'b0001110000111011100001111111111111111111111111111111111111110000,
    64'b0001110000111011100000000000000000000000000000000000000111111000,
    64'b0001110000111011100000000000000000000000000000000000000011111000,
    64'b0001110000111011100000000000000000000000000000000000000001111000,
    64'b0001110000111011111111111111111111111111111111111110000000111000,
    64'b0001110000111011111111111111111111111111111111111111100000111000,
    64'b0001110000111011111111111111111111111111111111111111110000111000,
    64'b0001110000111000000000000000000000000000000000001111110000111000,
    64'b0001110000111011111111111111111111111111111111111111100000111000,
    64'b0001110000111011111111111111111111111111111111111111100000111000,
    64'b0001110000111011111111111111111111111111111111111110000001111000,
    64'b0001110000111011100000000000000000000000000000000000000001111000,
    64'b0001110000111011100000000000000000000000000000000000000011111000,
    64'b0001110000111011100000000000000000000000000000000000000111110000,
    64'b0001110000111011100000000000000000000000000000000000011111110000,
    64'b0001110000111011100001111111111111111111111111111111111111100000,
    64'b0001110000111011100001111111111111111111111111111111111111100000,
    64'b0001110000111111100000000111111111111111111111111111111111110000,
    64'b0001110000111111100000000000000000000000000000000000000111110000,
    64'b0001110000111111110000000000000000000000000000000000000011110000,
    64'b0001110000011111111100000000000000000000000000000000000001110000,
    64'b0001110000011111111111100000000000000000000000000000000001110000,
    64'b0001111000001111111111111111111111111111111111111111100001110000,
    64'b0001111000000111111111111111111111111111111111111111100001110000,
    64'b0001111100000011111111111111111111111111111111111111100001110000,
    64'b0000111100000011111111111111111111111111111111111111100001110000,
    64'b0000111110000000111111111111111111111111111111111111100001110000,
    64'b0000011111000000000011111111111111111111111111111111100001110000,
    64'b0000011111100000000000000000000000000000000000000000000001110000,
    64'b0000001111111000000000000000000000000000000000000000000001110000,
    64'b0000000111111100000000000000000000000000000000000000000011110000,
    64'b0000000011111111100000000000000000000000000000000000000111110000,
    64'b0000000000111111111111111111111111111111111111111111111111110000,
    64'b0000000000011111111111111111111111111111111111111111111111100000,
    64'b0000000000000011111111111111111111111111111111111111111111000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000
};

logic [63:0] Emid_bitmap [0:63] = {
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000011111111111111111000000000000000000000000000,
    64'b0000000000000001111111111111111111111100000000000000000000000000,
    64'b0000000000000011111111111111111111111110000000000000000000000000,
    64'b0000000000001111111111111111111111111111000000000000000000000000,
    64'b0000000000011111111100000000000000001111000000000000000000000000,
    64'b0000000000111111000000000000000000001111000000000000000000000000,
    64'b0000000001111110000000000000000000001111000000000000000000000000,
    64'b0000000011111100000000000000000000001111000000000000000000000000,
    64'b0000000011111000000000000000000000001111010000000000000000000000,
    64'b0000000111110000000000000000000000001111000000000000000000000000,
    64'b0000001111100000000000000000000000001111000000000000000000000000,
    64'b0000001111000000000000011111111111111111000000000000000000000000,
    64'b0000001111000000000011111111111111111110000000000000000000000000,
    64'b0000001111000000000111111111111111111100000000000000000000000000,
    64'b0000001111000000000111111111111111111000000000000000000000000000,
    64'b0000001111000000011111110000000000000000000000000000000000000000,
    64'b0000001111000000011110000000000000000000000000000000000000000000,
    64'b0000001111000000011110000000000000000000000000000000000000000000,
    64'b0000001111000000011110000000000000000000000000000000000000000000,
    64'b0000001111000000011111111111111111111111111111111111111000000000,
    64'b0000001111000000011111111111111111111111111111111111111100000000,
    64'b0000001111000000011111111111111111111111111111111111111110000000,
    64'b0000001111000000000000000000000000000000000000000001111111000000,
    64'b0000001111000000000000000000000000000000000000000000011111000000,
    64'b0000001111000000000000000000000000000000000000000000001111000000,
    64'b0000001111000000000000000000000000000000000000000000001111000000,
    64'b0000001111000000000000000000000000000000000000000000011111000000,
    64'b0000001111000000000000000000000000000000000000000000011111000000,
    64'b0000001111000000000000000000000000000000000000000001111110000000,
    64'b0000001111000000011111111111111111111111111111111111111110000000,
    64'b0000001111000000011111111111111111111111111111111111111100000000,
    64'b0000001111000000011111111111111111111111111111111111111000000000,
    64'b0000001111000000011111111111111111111111111111111111100000000000,
    64'b0000001111000000011110000000000000000000000000000000000000000000,
    64'b0000001111000000011110000000000000000000000000000000000000000000,
    64'b0000001111000000011111111000000000000000000000000000000000000000,
    64'b0000001111000000011111111111111111111111111111111111111000000000,
    64'b0000001111000000001111111111111111111111111111111111111100000000,
    64'b0000001111100000000011111111111111111111111111111111111110000000,
    64'b0000001111100000000000011111111111111111111111111111111110000000,
    64'b0000000111110000000000000000000000000000000000000000011110000000,
    64'b0000000111111000000000000000000000000000000000000000011110000000,
    64'b0000000011111100000000000000000000000000000000000000011110000000,
    64'b0000000011111100000000000000000000000000000000000000011110000000,
    64'b0000000001111111000000000000000000000000000000000000011110000000,
    64'b0000000000111111111100000000000000000000000000000000011110000000,
    64'b0000000000011111111111111111111111111111111111111111111110000000,
    64'b0000000000000111111111111111111111111111111111111111111110000000,
    64'b0000000000000011111111111111111111111111111111111111111100000000,
    64'b0000000000000000011111111111111111111111111111111111111000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000
};

logic [63:0] Ein_bitmap [0:63] = {
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000011111111111111110000000000000000000000000000,
    64'b0000000000000000111111111111111111110000000000000000000000000000,
    64'b0000000000000001111111111111111111110000000000000000000000000000,
    64'b0000000000000011111111111111111111110000000000000000000000000000,
    64'b0000000000000111111111111111111111110000000000000000000000000000,
    64'b0000000000001111111111111111111111110000000000000000000000000000,
    64'b0000000000011111111111111111111111110000000000000000000000000000,
    64'b0000000000111111111111100000000000000000000000000000000000000000,
    64'b0000000000111111111100000000000000000000000000000000000000000000,
    64'b0000000000111111111000000000000000000000000000000000000000000000,
    64'b0000000000111111111000000000000000000000000000000000000000000000,
    64'b0000000000111111100000000000000000000000000000000000000000000000,
    64'b0000000000111111100000000000000000000000000000000000000000000000,
    64'b0000000000111111100000000000000000000000000000000000000000000000,
    64'b0000000000111111100000000000000000000000000000000000000000000000,
    64'b0000000000111111100000000000000000000000000000000000000000000000,
    64'b0000000000111111100000000000000000000000000000000000000000000000,
    64'b0000000000111111100000000000000000000000000000000000000000000000,
    64'b0000000000111111111111111111111111111111111111111110000000000000,
    64'b0000000000111111111111111111111111111111111111111111100000000000,
    64'b0000000000111111111111111111111111111111111111111111110000000000,
    64'b0000000000111111111111111111111111111111111111111111110000000000,
    64'b0000000000111111111111111111111111111111111111111111100000000000,
    64'b0000000000111111111111111111111111111111111111111111100000000000,
    64'b0000000000111111111111111111111111111111111111111110000000000000,
    64'b0000000000111111100000000000000000000000000000000000000000000000,
    64'b0000000000111111100000000000000000000000000000000000000000000000,
    64'b0000000000111111100000000000000000000000000000000000000000000000,
    64'b0000000000111111100000000000000000000000000000000000000000000000,
    64'b0000000000111111100000000000000000000000000000000000000000000000,
    64'b0000000000111111100000000000000000000000000000000000000000000000,
    64'b0000000000111111100000000000000000000000000000000000000000000000,
    64'b0000000000111111100000000000000000000000000000000000000000000000,
    64'b0000000000111111110000000000000000000000000000000000000000000000,
    64'b0000000000011111111100000000000000000000000000000000000000000000,
    64'b0000000000011111111111100000000000000000000000000000000000000000,
    64'b0000000000001111111111111111111111111111111111111111100000000000,
    64'b0000000000000111111111111111111111111111111111111111100000000000,
    64'b0000000000000011111111111111111111111111111111111111100000000000,
    64'b0000000000000011111111111111111111111111111111111111100000000000,
    64'b0000000000000000111111111111111111111111111111111111100000000000,
    64'b0000000000000000000011111111111111111111111111111111100000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000,
    64'b0000000000000000000000000000000000000000000000000000000000000000
};

    logic [31:0] Aout_bitmap32 [0:31] = {
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000011111111111111111111100000,
    32'b00000011111111111111111111100000,
    32'b00001100000000000000000000011000,
    32'b00001100000000000000000000011000,
    32'b00001100000011111111100000011000,
    32'b00001100000011111111100000011000,
    32'b00001100000011000001100000011000,
    32'b00001100000011000001100000011000,
    32'b00001100000011000001100000011000,
    32'b00001100000011000001100000011000,
    32'b00001100000011000001100000011000,
    32'b00001100000011000001100000011000,
    32'b00001100000011000001100000011000,
    32'b00001100000011111111100000011000,
    32'b00001100000011111111100000011000,
    32'b00001100000000000000000000011000,
    32'b00001100000000000000000000011000,
    32'b00001100000011111111100000011000,
    32'b00001100000011111111100000011000,
    32'b00001100000011000001100000011000,
    32'b00001100000011000001100000011000,
    32'b00001100000011000001100000011000,
    32'b00001100000011000001100000011000,
    32'b00001100000011000001100000011000,
    32'b00001100000011000001100000011000,
    32'b00001111111111000001111111111000,
    32'b00001111111111000001111111111000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000
};

logic [31:0] Ain_bitmap32 [0:31] = {
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000011111111111111111111100000,
    32'b00000011111111111111111111100000,
    32'b00000011111100000000011111100000,
    32'b00000011111100000000011111100000,
    32'b00000011111100000000011111100000,
    32'b00000011111100000000011111100000,
    32'b00000011111100000000011111100000,
    32'b00000011111100000000011111100000,
    32'b00000011111100000000011111100000,
    32'b00000011111100000000011111100000,
    32'b00000011111100000000011111100000,
    32'b00000011111100000000011111100000,
    32'b00000011111100000000011111100000,
    32'b00000011111111111111111111100000,
    32'b00000011111111111111111111100000,
    32'b00000011111100000000011111100000,
    32'b00000011111100000000011111100000,
    32'b00000011111100000000011111100000,
    32'b00000011111100000000011111100000,
    32'b00000011111100000000011111100000,
    32'b00000011111100000000011111100000,
    32'b00000011111100000000011111100000,
    32'b00000011111100000000011111100000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000
};

logic [31:0] Cout_bitmap32 [0:31] = {
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000111111111111111100000000,
    32'b00000000111111111111111100000000,
    32'b00000011000000000000000011000000,
    32'b00000011000000000000000011000000,
    32'b00000111000000000000000011100000,
    32'b00011000000111111111100000011000,
    32'b00011000000111111111100000011000,
    32'b00011000000110000001100000011000,
    32'b00011000000110000001111111111000,
    32'b00011000000110000001111111111000,
    32'b00011000000110000000000000000000,
    32'b00011000000110000000000000000000,
    32'b00011000000110000000000000000000,
    32'b00011000000110000000000000000000,
    32'b00011000000110000000000000000000,
    32'b00011000000110000000000000000000,
    32'b00011000000110000000000000000000,
    32'b00011000000110000000000000000000,
    32'b00011000000110000001111111111000,
    32'b00011000000110000001111111111000,
    32'b00011000000111111111100000011000,
    32'b00011000000111111111100000011000,
    32'b00011000000000000000000000011000,
    32'b00000111000000000000000011100000,
    32'b00000011000000000000000011000000,
    32'b00000000111111111111111100000000,
    32'b00000000111111111111111100000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000
};

logic [31:0] Cin_bitmap32 [0:31] = {
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000111111111111111100000000,
    32'b00000000111111111111111100000000,
    32'b00000000111111111111111100000000,
    32'b00000111111000000000011111100000,
    32'b00000111111000000000011111100000,
    32'b00000111111000000000011111100000,
    32'b00000111111000000000000000000000,
    32'b00000111111000000000000000000000,
    32'b00000111111000000000000000000000,
    32'b00000111111000000000000000000000,
    32'b00000111111000000000000000000000,
    32'b00000111111000000000000000000000,
    32'b00000111111000000000000000000000,
    32'b00000111111000000000000000000000,
    32'b00000111111000000000000000000000,
    32'b00000111111000000000000000000000,
    32'b00000111111000000000000000000000,
    32'b00000111111000000000000000000000,
    32'b00000111111000000000011111100000,
    32'b00000111111000000000011111100000,
    32'b00000111111111111111111111100000,
    32'b00000000111111111111111100000000,
    32'b00000000111111111111111100000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000
};


logic [31:0] Dout_bitmap32 [0:31] = {
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000111111111111111111000000000,
    32'b00000111111111111111111000000000,
    32'b00000110000000000000000110000000,
    32'b00000110000000000000000111000000,
    32'b00000110000011111000000000110000,
    32'b00000110000011111111000000110000,
    32'b00000110000011000011000000110000,
    32'b00000110000011000011000000110000,
    32'b00000110000011000011000000110000,
    32'b00000110000011000011000000110000,
    32'b00000110000011000011000000110000,
    32'b00000110000011000011000000110000,
    32'b00000110000011000011000000110000,
    32'b00000110000011000011000000110000,
    32'b00000110000011000011000000110000,
    32'b00000110000011000011000000110000,
    32'b00000110000011000011000000110000,
    32'b00000110000011000011000000110000,
    32'b00000110000011000011000000110000,
    32'b00000110000011111111000000110000,
    32'b00000110000011111111000000110000,
    32'b00000110000000000000000111000000,
    32'b00000110000000000000000110000000,
    32'b00000110000000000000000110000000,
    32'b00000111111111111111111000000000,
    32'b00000111111111111111111000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000
};

logic [31:0] Din_bitmap32 [0:31] = {
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000001111111111111111000000000,
    32'b00000001111111111111111000000000,
    32'b00000001111100000111111111000000,
    32'b00000001111100000000111111000000,
    32'b00000001111100000000111111000000,
    32'b00000001111100000000111111000000,
    32'b00000001111100000000111111000000,
    32'b00000001111100000000111111000000,
    32'b00000001111100000000111111000000,
    32'b00000001111100000000111111000000,
    32'b00000001111100000000111111000000,
    32'b00000001111100000000111111000000,
    32'b00000001111100000000111111000000,
    32'b00000001111100000000111111000000,
    32'b00000001111100000000111111000000,
    32'b00000001111100000000111111000000,
    32'b00000001111100000000111111000000,
    32'b00000001111100000000111111000000,
    32'b00000001111100000000111111000000,
    32'b00000001111111111111111000000000,
    32'b00000001111111111111111000000000,
    32'b00000001111111111111111000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000
};

logic [31:0] Eout_bitmap32 [0:31] = {
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00001111111111111111111111100000,
    32'b00001111111111111111111111100000,
    32'b00001100000000000000000001100000,
    32'b00001100000000000000000001100000,
    32'b00001100000111111111111111100000,
    32'b00001100000111111111111111100000,
    32'b00001100000110000000000000000000,
    32'b00001100000110000000000000000000,
    32'b00001100000110000000000000000000,
    32'b00001100000110000000000000000000,
    32'b00001100000111111111111110000000,
    32'b00001100000111111111111110000000,
    32'b00001100000000000000000110000000,
    32'b00001100000000000000000110000000,
    32'b00001100000111111111111110000000,
    32'b00001100000111111111111110000000,
    32'b00001100000110000000000000000000,
    32'b00001100000110000000000000000000,
    32'b00001100000110000000000000000000,
    32'b00001100000111111111111111100000,
    32'b00001100000111111111111111100000,
    32'b00001100000000000000000001100000,
    32'b00001100000000000000000001100000,
    32'b00001100000000000000000001100000,
    32'b00001111111111111111111111100000,
    32'b00001111111111111111111111100000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000
};


logic [31:0] Ein_bitmap32 [0:31] = {
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000011111111111111111110000000,
    32'b00000011111111111111111110000000,
    32'b00000011111000000000000000000000,
    32'b00000011111000000000000000000000,
    32'b00000011111000000000000000000000,
    32'b00000011111000000000000000000000,
    32'b00000011111000000000000000000000,
    32'b00000011111000000000000000000000,
    32'b00000011111000000000000000000000,
    32'b00000011111000000000000000000000,
    32'b00000011111111111111111000000000,
    32'b00000011111111111111111000000000,
    32'b00000011111000000000000000000000,
    32'b00000011111000000000000000000000,
    32'b00000011111000000000000000000000,
    32'b00000011111000000000000000000000,
    32'b00000011111000000000000000000000,
    32'b00000011111000000000000000000000,
    32'b00000011111000000000000000000000,
    32'b00000011111111111111111110000000,
    32'b00000011111111111111111110000000,
    32'b00000011111111111111111110000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000
};

logic [31:0] Fout_bitmap32 [0:31] = {
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000111111111111111111111110000,
    32'b00000111111111111111111111110000,
    32'b00000110000000000000000000110000,
    32'b00000110000000000000000000110000,
    32'b00000110000000000000000000110000,
    32'b00000110000011111111111111110000,
    32'b00000110000011111111111111110000,
    32'b00000110000011000000000000000000,
    32'b00000110000011000000000000000000,
    32'b00000110000011000000000000000000,
    32'b00000110000011111111111110000000,
    32'b00000110000011111111111110000000,
    32'b00000110000000000000000110000000,
    32'b00000110000000000000000110000000,
    32'b00000110000000000000000110000000,
    32'b00000110000011111111111110000000,
    32'b00000110000011111111111110000000,
    32'b00000110000011000000000000000000,
    32'b00000110000011000000000000000000,
    32'b00000110000011000000000000000000,
    32'b00000110000011000000000000000000,
    32'b00000110000011000000000000000000,
    32'b00000110000011000000000000000000,
    32'b00000110000011000000000000000000,
    32'b00000111111111000000000000000000,
    32'b00000111111111000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000
};

logic [31:0] Fin_bitmap32 [0:31] = {
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000001111111111111111111000000,
    32'b00000001111111111111111111000000,
    32'b00000001111111111111111111000000,
    32'b00000001111100000000000000000000,
    32'b00000001111100000000000000000000,
    32'b00000001111100000000000000000000,
    32'b00000001111100000000000000000000,
    32'b00000001111100000000000000000000,
    32'b00000001111100000000000000000000,
    32'b00000001111100000000000000000000,
    32'b00000001111111111111111000000000,
    32'b00000001111111111111111000000000,
    32'b00000001111111111111111000000000,
    32'b00000001111100000000000000000000,
    32'b00000001111100000000000000000000,
    32'b00000001111100000000000000000000,
    32'b00000001111100000000000000000000,
    32'b00000001111100000000000000000000,
    32'b00000001111100000000000000000000,
    32'b00000001111100000000000000000000,
    32'b00000001111100000000000000000000,
    32'b00000001111100000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000
};

logic [31:0] Lout_bitmap32 [0:31] = {
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00001111111111000000000000000000,
    32'b00001111111111000000000000000000,
    32'b00001100000011000000000000000000,
    32'b00001100000011000000000000000000,
    32'b00001100000011000000000000000000,
    32'b00001100000011000000000000000000,
    32'b00001100000011000000000000000000,
    32'b00001100000011000000000000000000,
    32'b00001100000011000000000000000000,
    32'b00001100000011000000000000000000,
    32'b00001100000011000000000000000000,
    32'b00001100000011000000000000000000,
    32'b00001100000011000000000000000000,
    32'b00001100000011000000000000000000,
    32'b00001100000011000000000000000000,
    32'b00001100000011000000000000000000,
    32'b00001100000011000000000000000000,
    32'b00001100000011000000000000000000,
    32'b00001100000011000000000000000000,
    32'b00001100000011000000000000000000,
    32'b00001100000011111111111111110000,
    32'b00001100000011111111111111110000,
    32'b00001100000000000000000000110000,
    32'b00001100000000000000000000110000,
    32'b00001111111111111111111111110000,
    32'b00001111111111111111111111110000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000
};

logic [31:0] Lin_bitmap32 [0:31] = {
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000011111100000000000000000000,
    32'b00000011111100000000000000000000,
    32'b00000011111100000000000000000000,
    32'b00000011111100000000000000000000,
    32'b00000011111100000000000000000000,
    32'b00000011111100000000000000000000,
    32'b00000011111100000000000000000000,
    32'b00000011111100000000000000000000,
    32'b00000011111100000000000000000000,
    32'b00000011111100000000000000000000,
    32'b00000011111100000000000000000000,
    32'b00000011111100000000000000000000,
    32'b00000011111100000000000000000000,
    32'b00000011111100000000000000000000,
    32'b00000011111100000000000000000000,
    32'b00000011111100000000000000000000,
    32'b00000011111100000000000000000000,
    32'b00000011111100000000000000000000,
    32'b00000011111100000000000000000000,
    32'b00000011111100000000000000000000,
    32'b00000011111111111111111111000000,
    32'b00000011111111111111111111000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000
};

logic [31:0] Nout_bitmap32 [0:31] = {
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000111111111111111111110000000,
    32'b00000111111111111111111110000000,
    32'b00000110000000000000000001100000,
    32'b00000110000000000000000001100000,
    32'b00000110000011111111000001100000,
    32'b00000110000011111111000001100000,
    32'b00000110000011000011000001100000,
    32'b00000110000011000011000001100000,
    32'b00000110000011000011000001100000,
    32'b00000110000011000011000001100000,
    32'b00000110000011000011000001100000,
    32'b00000110000011000011000001100000,
    32'b00000110000011000011000001100000,
    32'b00000110000011000011000001100000,
    32'b00000110000011000011000001100000,
    32'b00000110000011000011000001100000,
    32'b00000110000011000011000001100000,
    32'b00000110000011000011000001100000,
    32'b00000110000011000011000001100000,
    32'b00000110000011000011000001100000,
    32'b00000110000011000011000001100000,
    32'b00000110000011000011000001100000,
    32'b00000110000011000011000001100000,
    32'b00000110000011000011000001100000,
    32'b00000111111111000011111111100000,
    32'b00000111111111000011111111100000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000
};

logic [31:0] Nin_bitmap32 [0:31] = {
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000001111111111111111110000000,
    32'b00000001111111111111111110000000,
    32'b00000001111100000000111110000000,
    32'b00000001111100000000111110000000,
    32'b00000001111100000000111110000000,
    32'b00000001111100000000111110000000,
    32'b00000001111100000000111110000000,
    32'b00000001111100000000111110000000,
    32'b00000001111100000000111110000000,
    32'b00000001111100000000111110000000,
    32'b00000001111100000000111110000000,
    32'b00000001111100000000111110000000,
    32'b00000001111100000000111110000000,
    32'b00000001111100000000111110000000,
    32'b00000001111100000000111110000000,
    32'b00000001111100000000111110000000,
    32'b00000001111100000000111110000000,
    32'b00000001111100000000111110000000,
    32'b00000001111100000000111110000000,
    32'b00000001111100000000111110000000,
    32'b00000001111100000000111110000000,
    32'b00000001111100000000111110000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000
};

logic [31:0] Oout_bitmap32 [0:31] = {
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000001111111111111000000000,
    32'b00000000001111111111111000000000,
    32'b00000000110000000000000110000000,
    32'b00000001110000000000000111000000,
    32'b00000110000001111111000000110000,
    32'b00000110000001111111000000110000,
    32'b00000110000001100011000000110000,
    32'b00000110000001100011000000110000,
    32'b00000110000001100011000000110000,
    32'b00000110000001100011000000110000,
    32'b00000110000001100011000000110000,
    32'b00000110000001100011000000110000,
    32'b00000110000001100011000000110000,
    32'b00000110000001100011000000110000,
    32'b00000110000001100011000000110000,
    32'b00000110000001100011000000110000,
    32'b00000110000001100011000000110000,
    32'b00000110000001100011000000110000,
    32'b00000110000001100011000000110000,
    32'b00000110000001100011000000110000,
    32'b00000110000001111111000000110000,
    32'b00000110000001111111000000110000,
    32'b00000001110000000000000111000000,
    32'b00000000110000000000000110000000,
    32'b00000000001111111111111000000000,
    32'b00000000001111111111111000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000
};

logic [31:0] Oin_bitmap32 [0:31] = {
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000001111111111111000000000,
    32'b00000000001111111111111000000000,
    32'b00000001111110000000111111000000,
    32'b00000001111110000000111111000000,
    32'b00000001111110000000111111000000,
    32'b00000001111110000000111111000000,
    32'b00000001111110000000111111000000,
    32'b00000001111110000000111111000000,
    32'b00000001111110000000111111000000,
    32'b00000001111110000000111111000000,
    32'b00000001111110000000111111000000,
    32'b00000001111110000000111111000000,
    32'b00000001111110000000111111000000,
    32'b00000001111110000000111111000000,
    32'b00000001111110000000111111000000,
    32'b00000001111110000000111111000000,
    32'b00000001111110000000111111000000,
    32'b00000001111110000000111111000000,
    32'b00000001111110000000111111000000,
    32'b00000001111110000000111111000000,
    32'b00000000001111111111111000000000,
    32'b00000000001111111111111000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000
};

logic [31:0] Pout_bitmap32 [0:31] = {
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000001111111111111111110000000,
    32'b00000001111111111111111110000000,
    32'b00000110000000000000000001100000,
    32'b00000110000000000000000001100000,
    32'b00000110000011111111000001100000,
    32'b00000110000011111111000001100000,
    32'b00000110000011000011000001100000,
    32'b00000110000011000011000001100000,
    32'b00000110000011000011000001100000,
    32'b00000110000011000011000001100000,
    32'b00000110000011000011000001100000,
    32'b00000110000011000011000001100000,
    32'b00000110000011111111000001100000,
    32'b00000110000011111111000001100000,
    32'b00000110000000000000000001100000,
    32'b00000110000000000000000001100000,
    32'b00000110000011111111111110000000,
    32'b00000110000011111111111110000000,
    32'b00000110000011000000000000000000,
    32'b00000110000011000000000000000000,
    32'b00000110000011000000000000000000,
    32'b00000110000011000000000000000000,
    32'b00000110000011000000000000000000,
    32'b00000110000011000000000000000000,
    32'b00000111111111000000000000000000,
    32'b00000111111111000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000
};

logic [31:0] Pin_bitmap32 [0:31] = {
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000001111111111111111110000000,
    32'b00000001111111111111111110000000,
    32'b00000001111100000000111110000000,
    32'b00000001111100000000111110000000,
    32'b00000001111100000000111110000000,
    32'b00000001111100000000111110000000,
    32'b00000001111100000000111110000000,
    32'b00000001111100000000111110000000,
    32'b00000001111100000000111110000000,
    32'b00000001111100000000111110000000,
    32'b00000001111100000000111110000000,
    32'b00000001111100000000111110000000,
    32'b00000001111111111111111110000000,
    32'b00000001111111111111111110000000,
    32'b00000001111100000000000000000000,
    32'b00000001111100000000000000000000,
    32'b00000001111100000000000000000000,
    32'b00000001111100000000000000000000,
    32'b00000001111100000000000000000000,
    32'b00000001111100000000000000000000,
    32'b00000001111100000000000000000000,
    32'b00000001111100000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000
};

logic [31:0] Rout_bitmap32 [0:31] = {
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000001111111111111111100000000,
    32'b00000001111111111111111100000000,
    32'b00000110000000000000000011000000,
    32'b00000110000000000000000011000000,
    32'b00000110000000000000000011000000,
    32'b00000110000011111110000011000000,
    32'b00000110000011111110000011000000,
    32'b00000110000011000110000011000000,
    32'b00000110000011000110000011000000,
    32'b00000110000011000110000011000000,
    32'b00000110000011000110000011000000,
    32'b00000110000011000110000011000000,
    32'b00000110000011111110000011000000,
    32'b00000110000011111110000011000000,
    32'b00000110000000000000001100000000,
    32'b00000110000000000000001100000000,
    32'b00000110000000000000001100000000,
    32'b00000110000011111110000011000000,
    32'b00000110000011111110000011000000,
    32'b00000110000011000110000011000000,
    32'b00000110000011000110000011000000,
    32'b00000110000011000110000011000000,
    32'b00000110000011000110000011000000,
    32'b00000110000011000110000011000000,
    32'b00000111111111000111111111000000,
    32'b00000111111111000111111111000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000
};

logic [31:0] Rin_bitmap32 [0:31] = {
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000001111111111111111100000000,
    32'b00000001111111111111111100000000,
    32'b00000001111111111111111100000000,
    32'b00000001111100000001111100000000,
    32'b00000001111100000001111100000000,
    32'b00000001111100000001111100000000,
    32'b00000001111100000001111100000000,
    32'b00000001111100000001111100000000,
    32'b00000001111100000001111100000000,
    32'b00000001111100000001111100000000,
    32'b00000001111100000001111100000000,
    32'b00000001111100000001111100000000,
    32'b00000001111111111111110000000000,
    32'b00000001111111111111110000000000,
    32'b00000001111111111111110000000000,
    32'b00000001111100000001111100000000,
    32'b00000001111100000001111100000000,
    32'b00000001111100000001111100000000,
    32'b00000001111100000001111100000000,
    32'b00000001111100000001111100000000,
    32'b00000001111100000001111100000000,
    32'b00000001111100000001111100000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000
};

logic [31:0] Sout_bitmap32 [0:31] = {
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000011111111111111111000000,
    32'b00000000011111111111111111000000,
    32'b00000001100000000000000000110000,
    32'b00000001100000000000000000110000,
    32'b00000011100000000000000000110000,
    32'b00001100000011111111111111110000,
    32'b00001100000011111111111111110000,
    32'b00001100000011100000000000000000,
    32'b00001100000011100000000000000000,
    32'b00001100000011100000000000000000,
    32'b00001100000011111111111000000000,
    32'b00001100000011111111111000000000,
    32'b00000011100000000000000110000000,
    32'b00000001100000000000000111000000,
    32'b00000000011111111111000000110000,
    32'b00000000011111111111000000110000,
    32'b00000000000000000011000000110000,
    32'b00000000000000000011000000110000,
    32'b00000000000000000011000000110000,
    32'b00001111111111111111000000110000,
    32'b00001111111111111111000000110000,
    32'b00001100000000000000000111000000,
    32'b00001100000000000000000110000000,
    32'b00001100000000000000000110000000,
    32'b00000011111111111111111000000000,
    32'b00000011111111111111111000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000
};

logic [31:0] Sin_bitmap32 [0:31] = {
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000011111111111111111000000,
    32'b00000000011111111111111111000000,
    32'b00000000011111111111111111000000,
    32'b00000011111100000000000000000000,
    32'b00000011111100000000000000000000,
    32'b00000011111100000000000000000000,
    32'b00000011111100000000000000000000,
    32'b00000011111100000000000000000000,
    32'b00000011111100000000000000000000,
    32'b00000011111100000000000000000000,
    32'b00000011111111111111111000000000,
    32'b00000000011111111111111000000000,
    32'b00000000000000000000111111000000,
    32'b00000000000000000000111111000000,
    32'b00000000000000000000111111000000,
    32'b00000000000000000000111111000000,
    32'b00000000000000000000111111000000,
    32'b00000000000000000000111111000000,
    32'b00000000000000000000111111000000,
    32'b00000011111111111111111000000000,
    32'b00000011111111111111111000000000,
    32'b00000011111111111111111000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000
};

logic [31:0] Tout_bitmap32 [0:31] = {
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00001111111111111111111111111000,
    32'b00001111111111111111111111111000,
    32'b00001100000000000000000000011000,
    32'b00001100000000000000000000011000,
    32'b00001111111111000001111111111000,
    32'b00001111111111000001111111111000,
    32'b00000000000011000001100000000000,
    32'b00000000000011000001100000000000,
    32'b00000000000011000001100000000000,
    32'b00000000000011000001100000000000,
    32'b00000000000011000001100000000000,
    32'b00000000000011000001100000000000,
    32'b00000000000011000001100000000000,
    32'b00000000000011000001100000000000,
    32'b00000000000011000001100000000000,
    32'b00000000000011000001100000000000,
    32'b00000000000011000001100000000000,
    32'b00000000000011000001100000000000,
    32'b00000000000011000001100000000000,
    32'b00000000000011000001100000000000,
    32'b00000000000011000001100000000000,
    32'b00000000000011000001100000000000,
    32'b00000000000011000001100000000000,
    32'b00000000000011000001100000000000,
    32'b00000000000011111111100000000000,
    32'b00000000000011111111100000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000
};

logic [31:0] Tin_bitmap32 [0:31] = {
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000011111111111111111111100000,
    32'b00000011111111111111111111100000,
    32'b00000000000000111110000000000000,
    32'b00000000000000111110000000000000,
    32'b00000000000000111110000000000000,
    32'b00000000000000111110000000000000,
    32'b00000000000000111110000000000000,
    32'b00000000000000111110000000000000,
    32'b00000000000000111110000000000000,
    32'b00000000000000111110000000000000,
    32'b00000000000000111110000000000000,
    32'b00000000000000111110000000000000,
    32'b00000000000000111110000000000000,
    32'b00000000000000111110000000000000,
    32'b00000000000000111110000000000000,
    32'b00000000000000111110000000000000,
    32'b00000000000000111110000000000000,
    32'b00000000000000111110000000000000,
    32'b00000000000000111110000000000000,
    32'b00000000000000111110000000000000,
    32'b00000000000000111110000000000000,
    32'b00000000000000111110000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000
};

logic [31:0] Uout_bitmap32 [0:31] = {
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000111111111000011111111100000,
    32'b00000111111111000011111111100000,
    32'b00000110000000000000000001100000,
    32'b00000110000011000011000001100000,
    32'b00000110000011000011000001100000,
    32'b00000110000011000011000001100000,
    32'b00000110000011000011000001100000,
    32'b00000110000011000011000001100000,
    32'b00000110000011000011000001100000,
    32'b00000110000011000011000001100000,
    32'b00000110000011000011000001100000,
    32'b00000110000011000011000001100000,
    32'b00000110000011000011000001100000,
    32'b00000110000011000011000001100000,
    32'b00000110000011000011000001100000,
    32'b00000110000011000011000001100000,
    32'b00000110000011000011000001100000,
    32'b00000110000011000011000001100000,
    32'b00000110000011000011000001100000,
    32'b00000110000011111111000001100000,
    32'b00000110000011111111000001100000,
    32'b00000001110000000000000111000000,
    32'b00000000110000000000000110000000,
    32'b00000000110000000000000110000000,
    32'b00000000001111111111111000000000,
    32'b00000000001111111111111000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000
};

logic [31:0] Uin_bitmap32 [0:31] = {
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000001111100000000111110000000,
    32'b00000001111100000000111110000000,
    32'b00000001111100000000111110000000,
    32'b00000001111100000000111110000000,
    32'b00000001111100000000111110000000,
    32'b00000001111100000000111110000000,
    32'b00000001111100000000111110000000,
    32'b00000001111100000000111110000000,
    32'b00000001111100000000111110000000,
    32'b00000001111100000000111110000000,
    32'b00000001111100000000111110000000,
    32'b00000001111100000000111110000000,
    32'b00000001111100000000111110000000,
    32'b00000001111100000000111110000000,
    32'b00000001111100000000111110000000,
    32'b00000001111100000000111110000000,
    32'b00000001111100000000111110000000,
    32'b00000001111100000000111110000000,
    32'b00000001111100000000111110000000,
    32'b00000000001111111111111000000000,
    32'b00000000001111111111111000000000,
    32'b00000000001111111111111000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000
};

logic [31:0] Vout_bitmap32 [0:31] = {
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000001111111100001111111110000,
    32'b00000011111111100001111111110000,
    32'b00000110000001100001100000110000,
    32'b00000110000001100001100000110000,
    32'b00000110000001100001100000110000,
    32'b00000110000001100001100000110000,
    32'b00000110000001100001100000110000,
    32'b00000110000001100001100000110000,
    32'b00000110000001100001100000110000,
    32'b00000110000001100001100000110000,
    32'b00000110000001100001100000110000,
    32'b00000110000001100001100000110000,
    32'b00000110000001100001100000110000,
    32'b00000110000001100001100000110000,
    32'b00000110000001100001100000110000,
    32'b00000110000001100001100000110000,
    32'b00000110000001100001100000110000,
    32'b00000110000001100001100000110000,
    32'b00000110000001100011100000110000,
    32'b00000110000001111100000011000000,
    32'b00000110000001111100000011000000,
    32'b00000110000000000000000011000000,
    32'b00000110000000000000011100000000,
    32'b00000110000000000000011000000000,
    32'b00000111111111111111100000000000,
    32'b00000111111111111111100000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000
};

logic [31:0] Vin_bitmap32 [0:31] = {
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000001111110000000011111000000,
    32'b00000001111110000000011111000000,
    32'b00000001111110000000011111000000,
    32'b00000001111110000000011111000000,
    32'b00000001111110000000011111000000,
    32'b00000001111110000000011111000000,
    32'b00000001111110000000011111000000,
    32'b00000001111110000000011111000000,
    32'b00000001111110000000011111000000,
    32'b00000001111110000000011111000000,
    32'b00000001111110000000011111000000,
    32'b00000001111110000000011111000000,
    32'b00000001111110000000011111000000,
    32'b00000001111110000000011111000000,
    32'b00000001111110000000011111000000,
    32'b00000001111110000000011111000000,
    32'b00000001111110000000011111000000,
    32'b00000001111110000011111100000000,
    32'b00000001111110000011111100000000,
    32'b00000001111111111111111100000000,
    32'b00000001111111111111100000000000,
    32'b00000001111111111111100000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000
};


// w1_outer 레이어 비트맵 (32×32)
logic [31:0] Bout_bitmap32 [0:31] = {
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00011111111111111111111110000000,
    32'b00011111111111111111111110000000,
    32'b00011000000000000000000001100000,
    32'b00011000000000000000000001100000,
    32'b00011000000000000000000000110000,
    32'b00011000000111111111000000110000,
    32'b00011000000111111111000000110000,
    32'b00011000000111000111000000110000,
    32'b00011000000111000111000000110000,
    32'b00011000000111000111000000110000,
    32'b00011000000111111111000000110000,
    32'b00011000000111111111000000110000,
    32'b00011000000000000000000011100000,
    32'b00011000000000000000000011100000,
    32'b00011000000111111111000000110000,
    32'b00011000000111111111000000110000,
    32'b00011000000111000111000000110000,
    32'b00011000000111000111000000110000,
    32'b00011000000111000111000000110000,
    32'b00011000000111111111000000110000,
    32'b00011000000111111111000000110000,
    32'b00011000000000000000000001100000,
    32'b00011000000000000000000001100000,
    32'b00011000000000000000000001100000,
    32'b00011111111111111111111110000000,
    32'b00011111111111111111111110000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000
};

// w2_border 레이어 비트맵 (32×32)
logic [31:0] Bin_bitmap32 [0:31] = {
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000111111111111111111110000000,
    32'b00000111111111111111111110000000,
    32'b00000111111111111111111111000000,
    32'b00000111111000000000111111000000,
    32'b00000111111000000000111111000000,
    32'b00000111111000000000111111000000,
    32'b00000111111000000000111111000000,
    32'b00000111111000000000111111000000,
    32'b00000111111000000000111111000000,
    32'b00000111111000000000111111000000,
    32'b00000111111111111111111100000000,
    32'b00000111111111111111111100000000,
    32'b00000111111000000000111111000000,
    32'b00000111111000000000111111000000,
    32'b00000111111000000000111111000000,
    32'b00000111111000000000111111000000,
    32'b00000111111000000000111111000000,
    32'b00000111111000000000111111000000,
    32'b00000111111000000000111111000000,
    32'b00000111111111111111111100000000,
    32'b00000111111111111111111100000000,
    32'b00000111111111111111111100000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000
};

// w1_outer 레이어 비트맵 (32×32)
logic [31:0] Wout_bitmap32 [0:31] = {
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b11111111100000000000000111111110,
    32'b11111111100000000000000111111110,
    32'b11000001100011111111000110000110,
    32'b11000001100011111111000110000110,
    32'b11000001100011000011000110000110,
    32'b11000001100011000011000110000110,
    32'b11000001100011000011000110000110,
    32'b11000001100011000011000110000110,
    32'b11000001100011000011000110000110,
    32'b11000001100011000011000110000110,
    32'b11000001100011000011000110000110,
    32'b11000001100011000011000110000110,
    32'b11000001100011000011000110000110,
    32'b11000001100011000011000110000110,
    32'b11000001100011000011000110000110,
    32'b11000001100011000011000110000110,
    32'b11000001100011000011000110000110,
    32'b11000001100011000011000110000110,
    32'b11000001111100000000111110000110,
    32'b11100001111100000000111110000110,
    32'b11100001111100000000111110000110,
    32'b00111000000000111100000000011000,
    32'b00111000000000111100000000011000,
    32'b00111000000000111100000000011000,
    32'b00000111111111000011111111100000,
    32'b00000111111111000011111111100000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000
};

// w2_border 레이어 비트맵 (32×32)
logic [31:0] Win_bitmap32 [0:31] = {
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00111110000000000000000001111000,
    32'b00111110000000000000000001111000,
    32'b00111110000000111100000001111000,
    32'b00111110000000111100000001111000,
    32'b00111110000000111100000001111000,
    32'b00111110000000111100000001111000,
    32'b00111110000000111100000001111000,
    32'b00111110000000111100000001111000,
    32'b00111110000000111100000001111000,
    32'b00111110000000111100000001111000,
    32'b00111110000000111100000001111000,
    32'b00111110000000111100000001111000,
    32'b00111110000000111100000001111000,
    32'b00111110000000111100000001111000,
    32'b00111110000000111100000001111000,
    32'b00111110000000111100000001111000,
    32'b00111110000011111111000001111000,
    32'b00011110000011111111000001111000,
    32'b00011110000011111111000001111000,
    32'b00000111111111000011111111100000,
    32'b00000111111111000011111111100000,
    32'b00000111111111000011111111100000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000
};

// w1_outer 레이어 비트맵 (32×32)
logic [31:0] Yout_bitmap32 [0:31] = {
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00011111111110000001111111111000,
    32'b00011111111110000001111111111000,
    32'b00011000000110000001100000011000,
    32'b00011000000110000001100000011000,
    32'b00011000000110000001100000011000,
    32'b00011000000110000001100000011000,
    32'b00011000000110000001100000011000,
    32'b00011000000110000001100000011000,
    32'b00011000000110000001100000011000,
    32'b00000111000110000001100011100000,
    32'b00000111000111111111100011100000,
    32'b00000111000111111111100011100000,
    32'b00000000111000000000011100000000,
    32'b00000000111000000000011100000000,
    32'b00000000000111000011100000000000,
    32'b00000000000011000011000000000000,
    32'b00000000000011000011000000000000,
    32'b00000000000011000011000000000000,
    32'b00000000000011000011000000000000,
    32'b00000000000011000011000000000000,
    32'b00000000000011000011000000000000,
    32'b00000000000011000011000000000000,
    32'b00000000000011000011000000000000,
    32'b00000000000011000011000000000000,
    32'b00000000000011111111000000000000,
    32'b00000000000011111111000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000
};

// w2_border 레이어 비트맵 (32×32)
logic [31:0] Yin_bitmap32 [0:31] = {
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000111111000000000011111100000,
    32'b00000111111000000000011111100000,
    32'b00000111111000000000011111100000,
    32'b00000111111000000000011111100000,
    32'b00000111111000000000011111100000,
    32'b00000111111000000000011111100000,
    32'b00000111111000000000011111100000,
    32'b00000000111000000000011100000000,
    32'b00000000111000000000011100000000,
    32'b00000000111000000000011100000000,
    32'b00000000000111111111100000000000,
    32'b00000000000111111111100000000000,
    32'b00000000000000111100000000000000,
    32'b00000000000000111100000000000000,
    32'b00000000000000111100000000000000,
    32'b00000000000000111100000000000000,
    32'b00000000000000111100000000000000,
    32'b00000000000000111100000000000000,
    32'b00000000000000111100000000000000,
    32'b00000000000000111100000000000000,
    32'b00000000000000111100000000000000,
    32'b00000000000000111100000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000
};    

logic [31:0] zeroout_bitmap32 [0:31] = {
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000111111111111111110000000,
    32'b00000000111111111111111110000000,
    32'b00000011000000000000000011000000,
    32'b00000011000000000000000011000000,
    32'b00000011000000000000000011000000,
    32'b00000011000001111110000011000000,
    32'b00000011000001111110000011000000,
    32'b00000011000001100110000011000000,
    32'b00000011000001100110000011000000,
    32'b00000011000001100110000011000000,
    32'b00000011000001100110000011000000,
    32'b00000011000001100110000011000000,
    32'b00000011000001100110000011000000,
    32'b00000011000001100110000011000000,
    32'b00000011000001100110000011000000,
    32'b00000011000001100110000011000000,
    32'b00000011000001100110000011000000,
    32'b00000011000001100110000011000000,
    32'b00000011000001100110000011000000,
    32'b00000011000001111110000011000000,
    32'b00000011000001111110000011000000,
    32'b00000011000000000000000011000000,
    32'b00000011000000000000000011000000,
    32'b00000011000000000000000011000000,
    32'b00000000111111111111111100000000,
    32'b00000000111111111111111100000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000
};

    logic [31:0] zeroin_bitmap32 [0:31] = {
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000111111111111111100000000,
    32'b00000000111111111111111100000000,
    32'b00000000111111111111111100000000,
    32'b00000000111100000000111100000000,
    32'b00000000111100000000111100000000,
    32'b00000000111100000000111100000000,
    32'b00000000111100000000111100000000,
    32'b00000000111100000000111100000000,
    32'b00000000111100000000111100000000,
    32'b00000000111100000000111100000000,
    32'b00000000111100000000111100000000,
    32'b00000000111100000000111100000000,
    32'b00000000111100000000111100000000,
    32'b00000000111100000000111100000000,
    32'b00000000111100000000111100000000,
    32'b00000000111100000000111100000000,
    32'b00000000111100000000111100000000,
    32'b00000000111100000000111100000000,
    32'b00000000111100000000111100000000,
    32'b00000000111111111111111100000000,
    32'b00000000111111111111111100000000,
    32'b00000000111111111111111100000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000
};

// w1_outer 레이어 비트맵 (32×32)
logic [31:0] Hout_bitmap32 [0:31] = {
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00011111111110000001111111111000,
    32'b00011111111110000001111111111000,
    32'b00011000000110000001100000011000,
    32'b00011000000110000001100000011000,
    32'b00011000000110000001100000011000,
    32'b00011000000110000001100000011000,
    32'b00011000000110000001100000011000,
    32'b00011000000110000001100000011000,
    32'b00011000000110000001100000011000,
    32'b00011000000111111111100000011000,
    32'b00011000000111111111100000011000,
    32'b00011000000000000000000000011000,
    32'b00011000000000000000000000011000,
    32'b00011000000000000000000000011000,
    32'b00011000000111111111100000011000,
    32'b00011000000111111111100000011000,
    32'b00011000000110000001100000011000,
    32'b00011000000110000001100000011000,
    32'b00011000000110000001100000011000,
    32'b00011000000110000001100000011000,
    32'b00011000000110000001100000011000,
    32'b00011000000110000001100000011000,
    32'b00011000000110000001100000011000,
    32'b00011000000110000001100000011000,
    32'b00011111111110000001111111111000,
    32'b00011111111110000001111111111000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000
};

// w2_border 레이어 비트맵 (32×32)
logic [31:0] Hin_bitmap32 [0:31] = {
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000111111000000000011111100000,
    32'b00000111111000000000011111100000,
    32'b00000111111000000000011111100000,
    32'b00000111111000000000011111100000,
    32'b00000111111000000000011111100000,
    32'b00000111111000000000011111100000,
    32'b00000111111000000000011111100000,
    32'b00000111111000000000011111100000,
    32'b00000111111000000000011111100000,
    32'b00000111111111111111111111100000,
    32'b00000111111111111111111111100000,
    32'b00000111111111111111111111100000,
    32'b00000111111000000000011111100000,
    32'b00000111111000000000011111100000,
    32'b00000111111000000000011111100000,
    32'b00000111111000000000011111100000,
    32'b00000111111000000000011111100000,
    32'b00000111111000000000011111100000,
    32'b00000111111000000000011111100000,
    32'b00000111111000000000011111100000,
    32'b00000111111000000000011111100000,
    32'b00000111111000000000011111100000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000100,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000
};

// w1_outer 레이어 비트맵 (32×32)
logic [31:0] Iout_bitmap32 [0:31] = {
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00011111111111111111111111111000,
    32'b00011111111111111111111111111000,
    32'b00011000000000000000000000011000,
    32'b00011000000000000000000000011000,
    32'b00011000000000000000000000011000,
    32'b00011111111100000000111111111000,
    32'b00011111111100000000111111111000,
    32'b00000000001100000000110000000000,
    32'b00000000001100000000110000000000,
    32'b00000000001100000000110000000000,
    32'b00000000001100000000110000000000,
    32'b00000000001100000000110000000000,
    32'b00000000001100000000110000000000,
    32'b00000000001100000000110000000000,
    32'b00000000001100000000110000000000,
    32'b00000000001100000000110000000000,
    32'b00000000001100000000110000000000,
    32'b00000000001100000000110000000000,
    32'b00000000001100000000110000000000,
    32'b00011111111110000000111111111000,
    32'b00011111111110000000111111111000,
    32'b00011000000000000000000000011000,
    32'b00011000000000000000000000011000,
    32'b00011000000000000000000000011000,
    32'b00011111111111111111111111111000,
    32'b00011111111111111111111111111000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000
};

// w2_border 레이어 비트맵 (32×32)
logic [31:0] Iin_bitmap32 [0:31] = {
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000111111111111111111111100000,
    32'b00000111111111111111111111100000,
    32'b00000111111111111111111111100000,
    32'b00000000000011111111000000000000,
    32'b00000000000011111111000000000000,
    32'b00000000000011111111000000000000,
    32'b00000000000011111111000000000000,
    32'b00000000000011111111000000000000,
    32'b00000000000011111111000000000000,
    32'b00000000000011111111000000000000,
    32'b00000000000011111111000000000000,
    32'b00000000000011111111000000000000,
    32'b00000000000011111111000000000000,
    32'b00000000000011111111000000000000,
    32'b00000000000011111111000000000000,
    32'b00000000000011111111000000000000,
    32'b00000000000011111111000000000000,
    32'b00000000000011111111000000000000,
    32'b00000000000011111111000000000000,
    32'b00000111111111111111111111100000,
    32'b00000111111111111111111111100000,
    32'b00000111111111111111111111100000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000
};

// w1_outer 레이어 비트맵 (32×32)
logic [31:0] Gout_bitmap32 [0:31] = {
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000001111111111111111110000000,
    32'b00000001111111111111111110000000,
    32'b00000110000000000000000110000000,
    32'b00000110000000000000000110000000,
    32'b00011000000000000000000110000000,
    32'b00011000001111111111111110000000,
    32'b00011000001111111111111110000000,
    32'b00011000001100000000000000000000,
    32'b00011000001100000000000000000000,
    32'b00011000001100000000000000000000,
    32'b00011000001100001111111111110000,
    32'b00011000001100001111111111110000,
    32'b00011000001100001100000000110000,
    32'b00011000001100001100000000110000,
    32'b00011000001100001111111000110000,
    32'b00011000001100001111111000110000,
    32'b00011000001100000000011000110000,
    32'b00011000001100000000011000110000,
    32'b00011000001100000000011000110000,
    32'b00011000001111111111111000110000,
    32'b00011000001111111111111000110000,
    32'b00000110000000000000000000110000,
    32'b00000110000000000000000000110000,
    32'b00000110000000000000000000110000,
    32'b00000001111111111111111111000000,
    32'b00000001111111111111111111000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000
};

// w2_border 레이어 비트맵 (32×32)
logic [31:0] Gin_bitmap32 [0:31] = {
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000001111111111111111000000000,
    32'b00000001111111111111111000000000,
    32'b00000111111111111111111000000000,
    32'b00000111110000000000000000000000,
    32'b00000111110000000000000000000000,
    32'b00000111110000000000000000000000,
    32'b00000111110000000000000000000000,
    32'b00000111110000000000000000000000,
    32'b00000111110000000000000000000000,
    32'b00000111110000000000000000000000,
    32'b00000111110000000011111111000000,
    32'b00000111110000000011111111000000,
    32'b00000111110000000000000111000000,
    32'b00000111110000000000000111000000,
    32'b00000111110000000000000111000000,
    32'b00000111110000000000000111000000,
    32'b00000111110000000000000111000000,
    32'b00000111110000000000000111000000,
    32'b00000111110000000000000111000000,
    32'b00000001111111111111111111000000,
    32'b00000001111111111111111111000000,
    32'b00000001111111111111111111000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000
};

logic [31:0] Mout_bitmap32 [0:31] = {
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00111111111111111111111111111100,
    32'b00111111111111111111111111111100,
    32'b00110000000000000000000000001100,
    32'b00110000000000000000000000001100,
    32'b00110000000000000000000000001100,
    32'b00110000111111000011111100001100,
    32'b00110000111111000011111100001100,
    32'b00110000110011000011001100001100,
    32'b00110000110011000011001100001100,
    32'b00110000110011000011001100001100,
    32'b00110000110011000011001100001100,
    32'b00110000110011000011001100001100,
    32'b00110000110011000011001100001100,
    32'b00110000110011000011001100001100,
    32'b00110000110011000011001100001100,
    32'b00110000110011000011001100001100,
    32'b00110000110011000011001100001100,
    32'b00010000110011000011001100001100,
    32'b00110000110011000011001100001100,
    32'b00110000110011000011001100001100,
    32'b01110000110011000011001100001100,
    32'b00110000110011000011001100001100,
    32'b00110000110011000011001100001100,
    32'b00110000110011000011001100001100,
    32'b00111111110011111111001111111100,
    32'b00111111110011111111001111111100,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000
};

// w2_border 레이어 비트맵 (32×32)
logic [31:0] Min_bitmap32 [0:31] = {
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00001111111111111111111111110000,
    32'b00001111111111111111111111110000,
    32'b00001111111111111111111111110000,
    32'b00001111000000111100000011110000,
    32'b00001111000000111100000011110000,
    32'b00001111000000111100000011110000,
    32'b00001111000000111100000011110000,
    32'b00001111000000111100000011110000,
    32'b00001111000000111100000011110000,
    32'b00001111000000111100000011110000,
    32'b00001111000000111100000011110000,
    32'b00001111000000111100000011110000,
    32'b00001111000000111100000011110000,
    32'b00001111000000111100000011110000,
    32'b00001111000000111100000011110000,
    32'b01001111000000111100000011110000,
    32'b00001111000000111100000011110000,
    32'b00001111000000111100000011110000,
    32'b00001111000000111100000011110000,
    32'b00001111000000111100000011110000,
    32'b00001111000000111100000011110000,
    32'b00001111000000111100000011110000,
    32'b00001111000000111100000011110000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000
};

    logic [31:0] oneout_bitmap32 [0:31] = {
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000011111111111111100000000000,
    32'b00000011111111111111100000000000,
    32'b00000011000000000001100000000000,
    32'b00000011000000000001100000000000,
    32'b00000011000000000001100000000000,
    32'b00000011111111000001100000000000,
    32'b00000011111111000001100000000000,
    32'b00000000000011000001100000000000,
    32'b00000000000011000001100000000000,
    32'b00000000000011000001100000000000,
    32'b00000000000011000001100000000000,
    32'b00000000000011000001100000000000,
    32'b00000000000011000001100000000000,
    32'b00000000000011000001100000000000,
    32'b00000000000011000001100000000000,
    32'b00000000000011000001100000000000,
    32'b00000000000011000001100000000000,
    32'b00000000000011000001100000000000,
    32'b00000000000011000001100000000000,
    32'b00000011111111000001111111000000,
    32'b00000011111111000001111111000000,
    32'b00000011000000000000000011000000,
    32'b00000011000000000000000011000000,
    32'b00000011000000000000000011000000,
    32'b00000011111111111111111111000000,
    32'b00000011111111111111111111000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000
};

    logic [31:0] onein_bitmap32 [0:31] = {
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000111111111110000000000000,
    32'b00000000111111111110000000000000,
    32'b00000000111111111110000000000000,
    32'b00000000000000111110000000000000,
    32'b00000000000000111110000000000000,
    32'b00000000000000111110000000000000,
    32'b00000000000000111110000000000000,
    32'b00000000000000111110000000000000,
    32'b00000000000000111110000000000000,
    32'b00000000000000111110000000000000,
    32'b00000000000000111110000000000000,
    32'b00000000000000111110000000000000,
    32'b00000000000000111110000000000000,
    32'b00000000000000111110000000000000,
    32'b00000000000000111110000000000000,
    32'b00000000000000111110000000000000,
    32'b00000000000000111110000000000000,
    32'b00000000000000111110000000000000,
    32'b00000000000000111110000000000000,
    32'b00000000111111111111111100000000,
    32'b00000000111111111111111100000000,
    32'b00000000111111111111111100000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000
};

logic [31:0] twoout_bitmap32 [0:31] = {
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000001111111111111111000000000,
    32'b00000001111111111111111000000000,
    32'b00000110000000000000000110000000,
    32'b00000110000000000000000110000000,
    32'b00000110000000000000000001100000,
    32'b00000111111111111110000001100000,
    32'b00000111111111111110000001100000,
    32'b00000000000000000110000001100000,
    32'b00000000000000000110000001100000,
    32'b00000000000000000110000001100000,
    32'b00000000011111111110000001100000,
    32'b00000000011111111110000001100000,
    32'b00000001100000000000000110000000,
    32'b00000001100000000000000110000000,
    32'b00000001100000000000000110000000,
    32'b00000110000011111111111000000000,
    32'b00000110000011111111111000000000,
    32'b00000110000011000000000000000000,
    32'b00000110000011000000000000000000,
    32'b00000110000011100000000000000000,
    32'b00000110000011111111111111100000,
    32'b00000110000011111111111111100000,
    32'b00000110000000000000000001100000,
    32'b00000110000000000000000001100000,
    32'b00000110000000000000000001100000,
    32'b00000111111111111111111111100000,
    32'b00000111111111111111111111100000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000
};

logic [31:0] twoin_bitmap32 [0:31] = {
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000001111111111111111000000000,
    32'b00000001111111111111111000000000,
    32'b00000001111111111111111110000000,
    32'b00000000000000000000111110000000,
    32'b00000000000000000000111110000000,
    32'b00000000000000000000111110000000,
    32'b00000000000000000000111110000000,
    32'b00000000000000000000111110000000,
    32'b00000000000000000000111110000000,
    32'b00000000000000000000111110000000,
    32'b00000000011111111111111000000000,
    32'b00000000011111111111111000000000,
    32'b00000000011111111111111000000000,
    32'b00000001111100000000000000000000,
    32'b00000001111100000000000000000000,
    32'b00000001111100000000000000000000,
    32'b00000001111100000000000000000000,
    32'b00000001111100000000000000000000,
    32'b00000001111100000000000000000000,
    32'b00000001111100000000000000000000,
    32'b00000001111111111111111110000000,
    32'b00000001111111111111111110000000,
    32'b00000001111111111111111110000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000
};

logic [31:0] threeout_bitmap32 [0:31] = {
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000011111111111111111110000000,
    32'b00000011111111111111111110000000,
    32'b00001100000000000000000001100000,
    32'b00001100000000000000000001100000,
    32'b00001100000000000000000000011000,
    32'b00001111111111111111000000011000,
    32'b00001111111111111111000000011000,
    32'b00000000000000000011000000011000,
    32'b00000000000000000011000000011000,
    32'b00000000011111111111000000011000,
    32'b00000000011111111111000000011000,
    32'b00000000011000000000000001100000,
    32'b00000000011000000000000001100000,
    32'b00000000011000000000000001100000,
    32'b00000000011000000000000001100000,
    32'b00000000011111111111000000011000,
    32'b00000000011111111111000000011000,
    32'b00000000000000000011000000011000,
    32'b00000000000000000011000000011000,
    32'b00001111111111111111000000011000,
    32'b00001111111111111111000000011000,
    32'b00001100000000000000000000011000,
    32'b00001100000000000000000001100000,
    32'b00001100000000000000000001100000,
    32'b00000011111111111111111110000000,
    32'b00000011111111111111111110000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000
};

logic [31:0] threein_bitmap32 [0:31] = {
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000011111111111111111110000000,
    32'b00000011111111111111111110000000,
    32'b00000011111111111111111111100000,
    32'b00000000000000000000111111100000,
    32'b00000000000000000000111111100000,
    32'b00000000000000000000111111100000,
    32'b00000000000000000000111111100000,
    32'b00000000000000000000111111100000,
    32'b00000000000000000000111111100000,
    32'b00000000000111111111111110000000,
    32'b00000000000111111111111110000000,
    32'b00000000000111111111111110000000,
    32'b00000000000111111111111110000000,
    32'b00000000000000000000011111100000,
    32'b00000000000000000000011111100000,
    32'b00000000000000000000011111100000,
    32'b00000000000000000000011111100000,
    32'b00000000000000000000011111100000,
    32'b00000000000000000000011111100000,
    32'b00000011111111111111111111100000,
    32'b00000011111111111111111100000000,
    32'b00000011111111111111111100000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000
};

logic [31:0] fourout_bitmap32 [0:31] = {
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00001111111111000111111111100000,
    32'b00001111111111000111111111100000,
    32'b00001100000011000110000001100000,
    32'b00001100000011000110000001100000,
    32'b00001100000011000110000001100000,
    32'b00001100000011000110000001100000,
    32'b00001100000011000110000001100000,
    32'b00001100000011000110000001100000,
    32'b00001100000011000110000001100000,
    32'b00001100000011111110000001100000,
    32'b00001100000011111110000001100000,
    32'b00001100000000000000000001100000,
    32'b00001100000000000000000001100000,
    32'b00001100000000000000000001100000,
    32'b00001100000000000000000001100000,
    32'b00001111111111111110000001100000,
    32'b00001111111111111110000001100000,
    32'b00000000000000000110000001100000,
    32'b00000000000000000110000001100000,
    32'b00000000000000000110000001100000,
    32'b00000000000000000110000001100000,
    32'b00000000000000000110000001100000,
    32'b00000000000000000110000001100000,
    32'b00000000000000000110000001100000,
    32'b00000000000000000111111111100000,
    32'b00000000000000000111111111100000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000
};

logic [31:0] fourin_bitmap32 [0:31] = {
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000011111100000001111110000000,
    32'b00000011111100000001111110000000,
    32'b00000011111100000001111110000000,
    32'b00000011111100000001111110000000,
    32'b00000011111100000001111110000000,
    32'b00000011111100000001111110000000,
    32'b00000011111100000001111110000000,
    32'b00000011111100000001111110000000,
    32'b00000011111100000001111110000000,
    32'b00000011111111111111111110000000,
    32'b00000011111111111111111110000000,
    32'b00000011111111111111111110000000,
    32'b00000011111111111111111110000000,
    32'b00000000000000000001111110000000,
    32'b00000000000000000001111110000000,
    32'b00000000000000000001111110000000,
    32'b00000000000000000001111110000000,
    32'b00000000000000000001111110000000,
    32'b00000000000000000001111110000000,
    32'b00000000000000000001111110000000,
    32'b00000000000000000001111110000000,
    32'b00000000000000000001111110000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000
};

    logic [31:0] fiveout_bitmap32 [0:31] = {
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000111111111111111111111100000,
    32'b00000111111111111111111111100000,
    32'b00000110000000000000000001100000,
    32'b00000110000000000000000001100000,
    32'b00000110000000000000000001100000,
    32'b00000110000011111111111111100000,
    32'b00000110000011111111111111100000,
    32'b00000110000011100000000000000000,
    32'b00000110000011100000000000000000,
    32'b00000110000011111111111000000000,
    32'b00000110000011111111111000000000,
    32'b00000001100000000000000110000000,
    32'b00000001100000000000000110000000,
    32'b00000001100000000000000110000000,
    32'b00000000011111111111000001100000,
    32'b00000000011111111111000001100000,
    32'b00000000000000000011000001100000,
    32'b00000000000000000011000001100000,
    32'b00000000000000000011000001100000,
    32'b00000111111111111111000001100000,
    32'b00000111111111111111000001100000,
    32'b00000110000000000000000110000000,
    32'b00000110000000000000000110000000,
    32'b00000110000000000000000110000000,
    32'b00000001111111111111111000000000,
    32'b00000001111111111111111000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000
};

    logic [31:0] fivein_bitmap32 [0:31] = {
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000001111111111111111110000000,
    32'b00000001111111111111111110000000,
    32'b00000001111111111111111110000000,
    32'b00000001111100000000000000000000,
    32'b00000001111100000000000000000000,
    32'b00000001111100000000000000000000,
    32'b00000001111100000000000000000000,
    32'b00000001111100000000000000000000,
    32'b00000001111100000000000000000000,
    32'b00000000011111111111111000000000,
    32'b00000000011111111111111000000000,
    32'b00000000011111111111111000000000,
    32'b00000000000000000000111110000000,
    32'b00000000000000000000111110000000,
    32'b00000000000000000000111110000000,
    32'b00000000000000000000111110000000,
    32'b00000000000000000000111110000000,
    32'b00000000000000000000111110000000,
    32'b00000000000000000000111110000000,
    32'b00000001111111111111111000000000,
    32'b00000001111111111111111000000000,
    32'b00000001111111111111111000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000
};

    logic [31:0] sixout_bitmap32 [0:31] = {
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000111111111111111111000000,
    32'b00000000111111111111111111000000,
    32'b00000011000000000000000011000000,
    32'b00000011000000000000000011000000,
    32'b00000011000000000000000011000000,
    32'b00001100000011111111111111000000,
    32'b00001100000011111111111111000000,
    32'b00001100000011100000000000000000,
    32'b00001100000011100000000000000000,
    32'b00001100000011111111111110000000,
    32'b00001100000011111111111110000000,
    32'b00001100000000000000000001100000,
    32'b00001100000000000000000001100000,
    32'b00001100000000000000000001100000,
    32'b00001100000011111111100000011000,
    32'b00001100000011111111100000011000,
    32'b00001100000011000001100000011000,
    32'b00001100000011000001100000011000,
    32'b00001100000011111111100000011000,
    32'b00001100000011111111100000011000,
    32'b00000011000000000000000001100000,
    32'b00000011000000000000000001100000,
    32'b00000011000000000000000001100000,
    32'b00000000111111111111111110000000,
    32'b00000000111111111111111110000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000
};

    logic [31:0] sixin_bitmap32 [0:31] = {
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000111111111111111100000000,
    32'b00000000111111111111111100000000,
    32'b00000000111111111111111100000000,
    32'b00000011111100000000000000000000,
    32'b00000011111100000000000000000000,
    32'b00000011111100000000000000000000,
    32'b00000011111100000000000000000000,
    32'b00000011111100000000000000000000,
    32'b00000011111100000000000000000000,
    32'b00000011111111111111111110000000,
    32'b00000011111111111111111110000000,
    32'b00000011111111111111111110000000,
    32'b00000011111100000000011111100000,
    32'b00000011111100000000011111100000,
    32'b00000011111100000000011111100000,
    32'b00000011111100000000011111100000,
    32'b00000011111100000000011111100000,
    32'b00000011111100000000011111100000,
    32'b00000000111111111111111110000000,
    32'b00000000111111111111111110000000,
    32'b00000000111111111111111110000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000
};

logic [31:0] sevenout_bitmap32 [0:31] = {
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00001111111111111111111110000000,
    32'b00001111111111111111111110000000,
    32'b00001100000000000000000110000000,
    32'b00001100000000000000000110000000,
    32'b00001100000000000000000110000000,
    32'b00001111111111111000000110000000,
    32'b00001111111111111000000110000000,
    32'b00000000000000011000011000000000,
    32'b00000000000000011000011000000000,
    32'b00000000000011111001100000000000,
    32'b00000000000011111001100000000000,
    32'b00000000001100000110000000000000,
    32'b00000000001100000110000000000000,
    32'b00000000001100001100000000000000,
    32'b00000000001100011000000000000000,
    32'b00000000001100011000000000000000,
    32'b00000000001100011000000000000000,
    32'b00000000001100011000000000000000,
    32'b00000000001100011000000000000000,
    32'b00000000001100011000000000000000,
    32'b00000000001100011000000000000000,
    32'b00000000001100011000000000000000,
    32'b00000000001100011000000000000000,
    32'b00000000001100011000000000000000,
    32'b00000000001111111000000000000000,
    32'b00000000001111111000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000
};

logic [31:0] sevenin_bitmap32 [0:31] = {
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000011111111111111111000000000,
    32'b00000011111111111111111000000000,
    32'b00000011111111111111111000000000,
    32'b00000000000000000111111000000000,
    32'b00000000000000000111111000000000,
    32'b00000000000000000111100000000000,
    32'b00000000000000000111100000000000,
    32'b00000000000000000110000000000000,
    32'b00000000000000000110000000000000,
    32'b00000000000011111000000000000000,
    32'b00000000000011111000000000000000,
    32'b00000000000011110000000000000000,
    32'b00000000000011100000000000000000,
    32'b00000000000011100000000000000000,
    32'b00000000000011100000000000000000,
    32'b00000000000011100000000000000000,
    32'b00000000000011100000000000000000,
    32'b00000000000011100000000000000000,
    32'b00000000000011100000000000000000,
    32'b00000000000011100000000000000000,
    32'b00000000000011100000000000000000,
    32'b00000000000011100000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000
};

logic [31:0] eightout_bitmap32 [0:31] = {
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000011111111111111100000000,
    32'b00000000011111111111111100000000,
    32'b00000011000000000000000011000000,
    32'b00000011000000000000000011000000,
    32'b00001100000011111111000000110000,
    32'b00001100000011111111000000110000,
    32'b00001100000011100111000000110000,
    32'b00001100000011100111000000110000,
    32'b00001100000011100111000000110000,
    32'b00001100000011111111000000110000,
    32'b00001100000011111111000000110000,
    32'b00001100000011111111000000110000,
    32'b00000011000000000000000011000000,
    32'b00000011000000000000000011000000,
    32'b00000011000000000000000011000000,
    32'b00001100000011111111000000110000,
    32'b00001100000011111111000000110000,
    32'b00001100000011100111000000110000,
    32'b00001100000011100111000000110000,
    32'b00001100000011100111000000110000,
    32'b00001100000011111111000000110000,
    32'b00001100000011111111000000110000,
    32'b00000011000000000000000011000000,
    32'b00000011000000000000000011000000,
    32'b00000000111111111111111100000000,
    32'b00000000111111111111111100000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000
};

logic [31:0] eightin_bitmap32 [0:31] = {
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000111111111111111100000000,
    32'b00000000111111111111111100000000,
    32'b00000011111100000000111111000000,
    32'b00000011111100000000111111000000,
    32'b00000011111100000000111111000000,
    32'b00000011111100000000111111000000,
    32'b00000011111100000000111111000000,
    32'b00000011111100000000111111000000,
    32'b00000011111100000000111111000000,
    32'b00000011111100000000111111000000,
    32'b00000000111111111111111100000000,
    32'b00000000111111111111111100000000,
    32'b00000000111111111111111100000000,
    32'b00000001111100000000111111000000,
    32'b00000001111100000000111111000000,
    32'b00000001111100000000111111000000,
    32'b00000001111100000000111111000000,
    32'b00000001111100000000111111000000,
    32'b00000001111100000000111111000000,
    32'b00000001111100000000111111000000,
    32'b00000000011111111111111100000000,
    32'b00000000011111111111111100000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000
};

logic [31:0] nineout_bitmap32 [0:31] = {
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000001111111111110000000000,
    32'b00000000001111111111110000000000,
    32'b00000000110000000000001100000000,
    32'b00000000110000000000001100000000,
    32'b00000011000011111110000011000000,
    32'b00000011000011111110000011000000,
    32'b00000011000011000110000011000000,
    32'b00000011000011000110000011000000,
    32'b00000011000011000110000011000000,
    32'b00000011000011000110000011000000,
    32'b00000011000011111110000011000000,
    32'b00000011000011111110000011000000,
    32'b00000000110000000000000011000000,
    32'b00000000110000000000000011000000,
    32'b00000000001111111110000011000000,
    32'b00000000001111111110000011000000,
    32'b00000000000000000110000011000000,
    32'b00000000000000000110000011000000,
    32'b00000000000000000110000011000000,
    32'b00000000000000000110000011000000,
    32'b00000000000000000110000011000000,
    32'b00000000000000000110000011000000,
    32'b00000000000000000110000011000000,
    32'b00000000000000000110000011000000,
    32'b00000000000000000111111111000000,
    32'b00000000000000000111111111000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000
};

logic [31:0] ninein_bitmap32 [0:31] = {
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000001111111111110000000000,
    32'b00000000001111111111110000000000,
    32'b00000000111100000001111100000000,
    32'b00000000111100000001111100000000,
    32'b00000000111100000001111100000000,
    32'b00000000111100000001111100000000,
    32'b00000000111100000001111100000000,
    32'b00000000111100000001111100000000,
    32'b00000000111100000001111100000000,
    32'b00000000111100000001111100000000,
    32'b00000000001111111111111100000000,
    32'b00000000001111111111111100000000,
    32'b00000000000000000001111100000000,
    32'b00000000000000000001111100000000,
    32'b00000000000000000001111100000000,
    32'b00000000000000000001111100000000,
    32'b00000000000000000001111100000000,
    32'b00000000000000000001111100000000,
    32'b00000000000000000001111100000000,
    32'b00000000000000000001111100000000,
    32'b00000000000000000001111100000000,
    32'b00000000000000000001111100000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000
};

    logic [31:0] ex_bitmapout_32 [0:31] = {
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000111111111100000000000,
    32'b00000000000111111111100000000000,
    32'b00000000000110000001100000000000,
    32'b00000000000110000001100000000000,
    32'b00000000000110000001100000000000,
    32'b00000000000110000001100000000000,
    32'b00000000000110000001100000000000,
    32'b00000000000110000001100000000000,
    32'b00000000000110000001100000000000,
    32'b00000000000110000001100000000000,
    32'b00000000000110000001100000000000,
    32'b00000000000110000001100000000000,
    32'b00000000000110000001100000000000,
    32'b00000000000110000001100000000000,
    32'b00000000000110000001100000000000,
    32'b00000000000111111111100000000000,
    32'b00000000000111111111100000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000111111111100000000000,
    32'b00000000000111111111100000000000,
    32'b00000000000110000001100000000000,
    32'b00000000000110000001100000000000,
    32'b00000000000110000001100000000000,
    32'b00000000000110000001100000000000,
    32'b00000000000111111111100000000000,
    32'b00000000000111111111100000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000
};

// w2_border 레이어 비트맵 (32×32)
logic [31:0] ex_bitmapin_32 [0:31] = {
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000001111110000000000000,
    32'b00000000000001111110000000000000,
    32'b00000000000001111110000000000000,
    32'b00000000000001111110000000000000,
    32'b00000000000001111110000000000000,
    32'b00000000000001111110000000000000,
    32'b00000000000001111110000000000000,
    32'b00000000000001111110000000000000,
    32'b00000000000001111110000000000000,
    32'b00000000000001111110000000000000,
    32'b00000000000001111110000000000000,
    32'b00000000000001111110000000000000,
    32'b00000000000001111110000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000001111110000000000000,
    32'b00000000000001111110000000000000,
    32'b00000000000001111110000000000000,
    32'b00000000000001111110000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000
};

logic [31:0] co_bitmapout_32 [0:31] = {
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000001111111111110000000000,
    32'b00000000001111111111110000000000,
    32'b00000000001100000000110000000000,
    32'b00000000001100000000110000000000,
    32'b00000000001100000000110000000000,
    32'b00000000001100000000110000000000,
    32'b00000000001100000000110000000000,
    32'b00000000001111111111110000000000,
    32'b00000000001111111111110000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000001111111111110000000000,
    32'b00000000001111111111110000000000,
    32'b00000000001100000000110000000000,
    32'b00000000001100000000110000000000,
    32'b00000000001100000000110000000000,
    32'b00000000001100000000110000000000,
    32'b00000000001100000000110000000000,
    32'b00000000001111111111110000000000,
    32'b00000000001111111111110000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000
};
logic [31:0] co_bitmapin_32 [0:31] = {
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000011111111000000000000,
    32'b00000000000011111111000000000000,
    32'b00000000000011111111000000000000,
    32'b00000000000011111111000000000000,
    32'b00000000000011111111000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000011111111000000000000,
    32'b00000000000011111111000000000000,
    32'b00000000000011111111000000000000,
    32'b00000000000011111111000000000000,
    32'b00000000000011111111000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000
};
logic [31:0] dashout_bitmap32 [0:31] = {
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00011111111111111111111111111000,
    32'b00011111111111111111111111111000,
    32'b00011000000000000000000000011000,
    32'b00011000000000000000000000011000,
    32'b00011000000000000000000000011000,
    32'b00011000000000000000000000011000,
    32'b00011111111111111111111111111000,
    32'b00011111111111111111111111111000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000
};

logic [31:0] dashin_bitmap32 [0:31] = {
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000111111111111111111111100000,
    32'b00000111111111111111111111100000,
    32'b00000111111111111111111111100000,
    32'b00000111111111111111111111100000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000,
    32'b00000000000000000000000000000000
};

logic [21:0] black [0:21] = {
22'b0000000000000000000000,
22'b0000000000000000000000,
22'b0000111000000001111000,
22'b0001000111111110000100,
22'b0001000000000000000100,
22'b0001000000000000000100,
22'b0001000000000000000100,
22'b0000100000000000001000,
22'b0000100000000000001000,
22'b0000100000000000001000,
22'b0000100000000000001000,
22'b0000100010010000001000,
22'b0000100010010000001000,
22'b0000010000000000111000,
22'b0000001000000000100000,
22'b0000110000000000011000,
22'b0000100000000000001000,
22'b0000100000000011001000,
22'b0000111000000011111000,
22'b0000001000100010000000,
22'b0000000111011110000000,
22'b0000000000000000000000
};
logic [21:0] white [0:21] = {
22'b0000000000000000000000,
22'b0000000000000000000000,
22'b0000000000000000000000,
22'b0000111000000001111000,
22'b0000111111111111111000,
22'b0000111100001111111000,
22'b0000110100001001111000,
22'b0000000100001000010000,
22'b0000000100001000000000,
22'b0000001011110010000000,
22'b0000010000000001100000,
22'b0000010000000001110000,
22'b0000010000000001110000,
22'b0000001000000011000000,
22'b0000000111111111000000,
22'b0000000111111100000000,
22'b0000010111111100110000,
22'b0000011000000000110000,
22'b0000000000000000000000,
22'b0000000000000000000000,
22'b0000000000000000000000,
22'b0000000000000000000000
};
logic [21:0] green [0:21] = {
22'b0000000000000000000000,
22'b0000000000000000000000,
22'b0000000000000000000000,
22'b0000000000000000000000,
22'b0000000000000000000000,
22'b0000000011110000000000,
22'b0000001011110110000000,
22'b0000011011110111100000,
22'b0000010000000001110000,
22'b0000000000000000010000,
22'b0000000000000000000000,
22'b0000000000000000000000,
22'b0000000000000000000000,
22'b0000000000000000000000,
22'b0000000000000000000000,
22'b0000000000000000000000,
22'b0000000000000000000000,
22'b0000000000000000000000,
22'b0000000111111100000000,
22'b0000000111011100000000,
22'b0000000000000000000000,
22'b0000000000000000000000
};
logic [21:0] lime [0:21] = {
22'b0000000000000000000000,
22'b0000000000000000000000,
22'b0000000000000000000000,
22'b0000000000000000000000,
22'b0000000000000000000000,
22'b0000000000000000000000,
22'b0000000000000000000000,
22'b0000000000000000000000,
22'b0000001011110110000000,
22'b0000010000000001100000,
22'b0000000000000000010000,
22'b0000000000000000000000,
22'b0000000000000000000000,
22'b0000000000000000000000,
22'b0000000000000000000000,
22'b0000000000000000000000,
22'b0000000000000000000000,
22'b0000000101110100000000,
22'b0000000000000000000000,
22'b0000000000000000000000,
22'b0000000000000000000000,
22'b0000000000000000000000
};
logic [21:0] skin [0:21] = {
22'b0000000000000000000000,
22'b0000000000000000000000,
22'b0000000000000000000000,
22'b0000000000000000000000,
22'b0000000000000000000000,
22'b0000000000000000000000,
22'b0000000000000000000000,
22'b0000000000000000000000,
22'b0000000000000000000000,
22'b0000000100001100000000,
22'b0000001111111110000000,
22'b0000001101101110000000,
22'b0000000001100010000000,
22'b0000000110011100000000,
22'b0000000000000000000000,
22'b0000001000000011100000,
22'b0000001000000011000000,
22'b0000000000000000000000,
22'b0000000000000000000000,
22'b0000000000000000000000,
22'b0000000000000000000000,
22'b0000000000000000000000
};
logic [21:0] pink [0:21] = {
22'b0000000000000000000000,
22'b0000000000000000000000,
22'b0000000000000000000000,
22'b0000000000000000000000,
22'b0000000000000000000000,
22'b0000000000000000000000,
22'b0000000000000000000000,
22'b0000000000000000000000,
22'b0000000000000000000000,
22'b0000000000000000000000,
22'b0000000000000000000000,
22'b0000000000000000000000,
22'b0000001100001100000000,
22'b0000000000000000000000,
22'b0000000000000000000000,
22'b0000000000000000000000,
22'b0000000000000000000000,
22'b0000000000000000000000,
22'b0000000000000000000000,
22'b0000000000000000000000,
22'b0000000000000000000000,
22'b0000000000000000000000
};
logic [21:0] yellow [0:21] = {
22'b0000000000000000000000,
22'b0000000000000000000000,
22'b0000000000000000000000,
22'b0000000000000000000000,
22'b0000000000000000000000,
22'b0000000000000000000000,
22'b0000000000000000000000,
22'b0000000000000000000000,
22'b0000000000000000000000,
22'b0000000000000000000000,
22'b0000000000000000000000,
22'b0000000000000000000000,
22'b0000000000000000000000,
22'b0000000001100000000000,
22'b0000000000000000000000,
22'b0000000000000000000000,
22'b0000000000000000000000,
22'b0000000010001000000000,
22'b0000000000000000000000,
22'b0000000000000000000000,
22'b0000000000000000000000,
22'b0000000000000000000000
};
//////////////////////////------------STATE---------------//////////////////////////////////////////////////////////////////////
    localparam IDLE = 0, SEL_LEVEL = 1, LEVEL0 = 2, LEVEL1_1 = 3, LEVEL1_2 = 4, LEVEL1_3 = 5,
    LEVEL2_1 = 6, LEVEL2_2 = 7, LEVEL2_3 = 8, WIN_LOSE = 9, WIN_DSIPLAY = 10, LOSE_DSIPLAY = 11, START = 12, GAME_DONE = 13, HOLD = 14, HOLD2 = 15,
    LEVEL3_1 = 16, LEVEL3_2 = 17, LEVEL3_3 = 18, END_DISPLAY = 19;
    logic [4:0] state, state_next;
//////////////////////////------------STATE---------------//////////////////////////////////////////////////////////////////////


//////////////////////////------------FONT LOCATION AND COLOR-----------//////////////////////////////////////////////////////////////////////
    logic [2:0] x_off, y_off; // x,y offset 글자 비트맵 통해서 1인 부분만 출력하기 위해
    logic [4:0] x_32, y_32;
    logic [5:0] x_64, y_64;
    logic w_mid, w_in, w_out, L_in, L_mid, L_out, font_in, font_out, R_in, Y_in, B_in, G_in, P_in, White_in, countcolor_in,
          cha_1, cha_2, cha_3, cha_4, cha_5, cha_6, cha_7; // 비트맵의의 1인 부분을 rgb 포트를 통해서 색깔 정함



    localparam RUNFORCOLOR_X = 100, RUNFORCOLOR_Y = 20, SPACE_3= 3, BIT31 = 31, SPACE_32=32;

//////////////////////////------------FONT LOCATION AND COLOR-----------//////////////////////////////////////////////////////////////////////


//////////////////////////------------ SCORE -----------//////////////////////////////////////////////////////////////////////
    logic zero_in, zero_out, one_in, one_out, two_in, two_out, three_in, three_out,
        four_in, four_out, five_in, five_out, six_in, six_out, seven_in, seven_out, eight_in, eight_out, nine_in, nine_out;
    logic [3:0] score, score_next;
    logic [3:0] high_score, high_score_next;
    logic give_done_ff1, give_done_ff2;
    logic start_ff1, start_ff2;
//////////////////////////------------ SCORE -----------//////////////////////////////////////////////////////////////////////


//////////////////////////------------FONT LOCATION AND COLOR-----------//////////////////////////////////////////////////////////////////////


//////////////////////////---------------COUNT-------------------//////////////////////////////////////////////////////////////////////
    logic [$clog2(25_000_000)-1:0]
        clk_counter, clk_counter_next, clk_counter_blink, clk_counter_blink_next, clk_counter_delay, clk_counter_delay_next, clk_counter_end, clk_counter_end_next;  // 25MHz 기준으로 1초 카운터

    logic hold_counter, hold_counter_next;
    // logic [3:0] countdown, countdown_next;  // 카운트다운 타이머
    logic [3:0] countdown_next, countdown_end, countdown_end_next;  // 카운트다운 타이머
    logic [5:0] blink_count, blink_count_next; // 0.2초 깜빡이기 위한 카운터
    logic [3:0] delay_count, delay_count_next;
    // logic [1:0] startcount, startcount_next;  // 시작 카운트
    logic [1:0] startcount_next;  // 시작 카운트
    logic [3:0] lvl_count, lvl_count_next;

    logic [$clog2(25_000_000)-1:0] frame_counter, frame_counter_next;
    logic [9:0] frame, frame_next;

    logic
        countdown_done_reg,
        countdown_done_next;  // 카운트다운 완료 신호,
    logic game_done_reg, game_done_next;  // 게임 완료 신호
    logic give_comparison_done_next;
    logic q_display_done, q_display_done_next;

    logic [3:0] led_next;

    logic end_reg, end_next;

    assign countdown_done = countdown_done_reg;
    assign slave_done = game_done_reg;
//////////////////////////---------------COUNT-------------------//////////////////////////////////////////////////////////////////////


//////////////////////////---------------ANIMATION-------------------//////////////////////////////////////////////////////////////////////
    logic [9:0] temp_x_coordinate, temp_x_coordinate_next;
    logic [9:0] temp_y_coordinate, temp_y_coordinate_next;

    // FRAME, 0.1sec
    localparam FRAMECOUNTER = 2_500_000; 

    //LETTER DEFAULT VALUE
    localparam LETTER_INTERVAL = 6;
    localparam WIDTH64 = 64;
    localparam WIDTH32 = 32;


    // WIN/LOSE LETTER
    localparam WL_DISPLAY_Y1 = 88, WL_DISPLAY_Y2 = 152;
    localparam W_X_COORDINATE = 196;
    localparam L_X_COORDINATE = 145;


    // LEVEL LETTER
    localparam LVL_X_COORDINATE = 0; 
    localparam LVL_Y_COORDINATE = 0; 

    // SCORE LETTER
    localparam SCORE_X_COORDINATE = 525;

//////////////////////////---------------ANIMATION-------------------//////////////////////////////////////////////////////////////////////



    always_ff @(posedge pclk, posedge reset) begin
        if (reset) begin
            state <= IDLE;  // 초기 상태
            clk_counter <= 0;  // 카운터 초기화
            clk_counter_blink <= 0; // 카운터 초기화화
            clk_counter_delay <= 0;
            clk_counter_end <= 0;
            countdown <= 5;  // 초 단위 초기화 
            startcount <= 3;  // 시작 카운트 초기화
            countdown_end <= 10;
            game_done_reg <= 1;  // 게임 완료 신호 초기화
            countdown_done_reg <= 0; // 카운트다운 완료 신호 초기화
            blink_count <= 0;   // 블링크 카운트 신호 초기화화
            delay_count <= 0;
            give_comparison_done <= 0;
            q_display_done <= 0;
            frame_counter <= 0;
            frame <= 0;
            temp_x_coordinate <= 0;
            temp_y_coordinate <= 0;
            score <= 0;
            high_score <= 0;
            test_led <= 0;
            // score
            score <= 0;
            lvl_count <= 0;
            end_reg <= 0;
        end else begin
            state <= state_next;  // 상태 업데이트
            countdown <= countdown_next;
            startcount <= startcount_next;  // 시작 카운트 업데이트
            clk_counter <= clk_counter_next;  // 카운터 증가
            clk_counter_blink <= clk_counter_blink_next;
            clk_counter_end <= clk_counter_end_next;
            game_done_reg <= game_done_next;  // 게임 완료 신호 업데이트
            countdown_done_reg <= countdown_done_next;
            blink_count <= blink_count_next;
            clk_counter_delay <= clk_counter_delay_next;
            delay_count <= delay_count_next;
            countdown_end <= countdown_end_next;
            give_comparison_done <= give_comparison_done_next;
            q_display_done <= q_display_done_next;
            frame_counter <= frame_counter_next;
            frame <= frame_next;
            temp_x_coordinate <= temp_x_coordinate_next;
            temp_y_coordinate <= temp_y_coordinate_next;
            score <= score_next;
            high_score <= high_score_next;
            test_led <= led_next;
            start_ff1 <= sw;
            start_ff2 <= start_ff1;
            give_done_ff1 <= give_done;
            give_done_ff2 <= give_done_ff1;
            lvl_count <= lvl_count_next;
            end_reg <= end_next;
        end
    end


    always_comb begin
        red_port = cam_r;  // 카메라 입력값
        green_port = cam_g;  // 카메라 입력값
        blue_port = cam_b;  // 카메라 입력값
        state_next = state;  // 상태 초기화
        clk_counter_next = clk_counter;
        clk_counter_blink_next = clk_counter_blink;
        clk_counter_delay_next = clk_counter_delay;
        clk_counter_end_next = clk_counter_end;
        countdown_next = countdown;  // 카운트다운 초기화
        blink_count_next = blink_count;
        countdown_end_next = countdown_end;
        startcount_next = startcount;  // 시작 카운트 초기화
        countdown_done_next = countdown_done_reg;  // 카운트다운 완료 신호 초기화
        game_done_next = game_done_reg;  // 게임 완료 신호 초기화
        delay_count_next = delay_count;
        hold_counter_next = hold_counter;
        give_comparison_done_next = give_comparison_done;
        q_display_done_next = q_display_done;
        frame_counter_next = frame_counter;
        frame_next = frame;
        temp_x_coordinate_next = temp_x_coordinate;
        temp_y_coordinate_next = temp_y_coordinate;
        // score
        score_next = score;
        high_score_next = high_score;
        led_next = test_led;
        lvl_count_next = lvl_count;
        end_next = end_reg;
        w_in = 0;
        w_mid = 0;   
        w_out = 0;
        L_in = 0;
        L_mid = 0;
        L_out = 0;
        font_in = 0;
        font_out = 0;
        R_in = 0;
        Y_in = 0;
        B_in = 0;
        G_in = 0;
        P_in = 0;
        White_in = 0;
        cha_1 = 0;
        cha_2 = 0;
        cha_3 = 0;
        cha_4 = 0;
        cha_5 = 0;
        cha_6 = 0;
        cha_7 = 0;
        countcolor_in = 0;

        bgm_enable = (state == IDLE || state == END_DISPLAY);              


        case (state)
        /************************************IDLE******************************************/
        /************************************IDLE******************************************/
        /************************************IDLE******************************************/
        /************************************IDLE******************************************/
        /************************************IDLE******************************************/
        /************************************IDLE******************************************/
        /************************************IDLE******************************************/
        /************************************IDLE******************************************/
        /************************************IDLE******************************************/
        /************************************IDLE******************************************/
            IDLE: // 게임 시작 전 로딩 화면
            begin
                countdown_done_next = 0;  // 카운트다운 완료 신호 초기화
                game_done_next = 1;  // 게임 완료 신호 초기화
                hold_counter_next = 0;
                give_comparison_done_next = 0;
                frame_next = 0;
                temp_x_coordinate_next = 0;
                temp_y_coordinate_next = 0;
                led_next = 4'b0111;
                score_next = 0;
                countdown_next = 5;
                startcount_next =3;
                countdown_end_next = 10;
                // 게임 제목 "Run For Color" 출력
                // RUNFORCOLOR_X = 100, RUNFORCOLOR_Y = 20, SPACE_3= 3, BIT31 = 31 SPACE_32=32;
                if (y_pixel >= RUNFORCOLOR_Y && y_pixel < RUNFORCOLOR_Y + SPACE_32 ) begin 
                    y_32 = y_pixel - RUNFORCOLOR_Y;

                    case (x_pixel) inside
                    [(RUNFORCOLOR_X):(RUNFORCOLOR_X + BIT31)] : begin //  100 ~ 131                  
                        x_32 = x_pixel - (RUNFORCOLOR_X);
                        font_out = Rout_bitmap32[y_32][31-x_32];
                        font_in = Rin_bitmap32[y_32][31-x_32];
                    end
                    [(RUNFORCOLOR_X + BIT31 + SPACE_3):(RUNFORCOLOR_X + 2*BIT31 + SPACE_3)] : begin //  134 ~ 165
                        x_32 = x_pixel - (RUNFORCOLOR_X+ BIT31 +SPACE_3);
                        font_out = Uout_bitmap32[y_32][31-x_32];
                        font_in = Uin_bitmap32[y_32][31-x_32];
                    end 
                    [(RUNFORCOLOR_X + 2*BIT31 + 2*SPACE_3):(RUNFORCOLOR_X + 3*BIT31 + 2*SPACE_3)] : begin // 168 ~ 199
                        x_32 = x_pixel - (RUNFORCOLOR_X + 2*BIT31 + 2*SPACE_3);
                        font_out = Nout_bitmap32[y_32][31-x_32];
                        font_in = Nin_bitmap32[y_32][31-x_32];
                    end
                    //space32
                    [(RUNFORCOLOR_X + 3*BIT31 + 3*SPACE_3 + SPACE_32):(RUNFORCOLOR_X + 4*BIT31 + 3*SPACE_3 + SPACE_32)] : begin // 168 ~ 199
                        x_32 = x_pixel - (RUNFORCOLOR_X + 3*BIT31 + 3*SPACE_3 + SPACE_32);
                        font_out = Fout_bitmap32[y_32][31-x_32];
                        font_in = Fin_bitmap32[y_32][31-x_32];
                    end
                    [(RUNFORCOLOR_X + 4*BIT31 + 4*SPACE_3 + SPACE_32):(RUNFORCOLOR_X + 5*BIT31 + 4*SPACE_3 + SPACE_32)] : begin // 168 ~ 199
                        x_32 = x_pixel - (RUNFORCOLOR_X + 4*BIT31 + 4*SPACE_3 + SPACE_32);
                        font_out = Oout_bitmap32[y_32][31-x_32];
                        font_in = Oin_bitmap32[y_32][31-x_32];
                    end
                    [(RUNFORCOLOR_X + 5*BIT31 + 5*SPACE_3 + SPACE_32):(RUNFORCOLOR_X + 6*BIT31 + 5*SPACE_3 + SPACE_32)] : begin // 168 ~ 199
                        x_32 = x_pixel - (RUNFORCOLOR_X + 5*BIT31 + 5*SPACE_3 + SPACE_32);
                        font_out = Rout_bitmap32[y_32][31-x_32];
                        font_in = Rin_bitmap32[y_32][31-x_32];
                    end
                    //space32
                    [(RUNFORCOLOR_X + 6*BIT31 + 6*SPACE_3 + 2*SPACE_32):(RUNFORCOLOR_X + 7*BIT31 + 6*SPACE_3 + 2*SPACE_32)] : begin // 168 ~ 199
                        x_32 = x_pixel - (RUNFORCOLOR_X + 6*BIT31 + 6*SPACE_3 + 2*SPACE_32);
                        font_out = Cout_bitmap32[y_32][31-x_32];
                        font_in = Cin_bitmap32[y_32][31-x_32];
                    end
                    [(RUNFORCOLOR_X + 7*BIT31 + 7*SPACE_3 + 2*SPACE_32):(RUNFORCOLOR_X + 8*BIT31 + 7*SPACE_3 + 2*SPACE_32)] : begin // 168 ~ 199
                        x_32 = x_pixel - (RUNFORCOLOR_X + 7*BIT31 + 7*SPACE_3 + 2*SPACE_32);
                        font_out = Oout_bitmap32[y_32][31-x_32];
                        font_in = Oin_bitmap32[y_32][31-x_32];
                    end
                    [(RUNFORCOLOR_X + 8*BIT31 + 8*SPACE_3 + 2*SPACE_32):(RUNFORCOLOR_X + 9*BIT31 + 8*SPACE_3 + 2*SPACE_32)] : begin // 168 ~ 199
                        x_32 = x_pixel - (RUNFORCOLOR_X + 8*BIT31 + 8*SPACE_3 + 2*SPACE_32);
                        font_out = Lout_bitmap32[y_32][31-x_32];
                        font_in = Lin_bitmap32[y_32][31-x_32];
                    end
                    [(RUNFORCOLOR_X + 9*BIT31 + 9*SPACE_3 + 2*SPACE_32):(RUNFORCOLOR_X + 10*BIT31 + 9*SPACE_3 + 2*SPACE_32)] : begin // 168 ~ 199
                        x_32 = x_pixel - (RUNFORCOLOR_X + 9*BIT31 + 9*SPACE_3 + 2*SPACE_32);
                        font_out = Oout_bitmap32[y_32][31-x_32];
                        font_in = Oin_bitmap32[y_32][31-x_32];
                    end
                    [(RUNFORCOLOR_X + 10*BIT31 + 10*SPACE_3 + 2*SPACE_32):(RUNFORCOLOR_X + 11*BIT31 + 10*SPACE_3 + 2*SPACE_32)] : begin // 168 ~ 199
                        x_32 = x_pixel - (RUNFORCOLOR_X + 10*BIT31 + 10*SPACE_3 + 2*SPACE_32);
                        font_out = Rout_bitmap32[y_32][31-x_32];
                        font_in = Rin_bitmap32[y_32][31-x_32];
                    end
                    endcase
                end else if (y_pixel >= 324 && y_pixel < 356 ) begin 
                    y_32 = y_pixel - 324;
                    case (x_pixel) inside
                    [100:131] : begin                  
                        x_32 = x_pixel - (100);
                        font_out = Hout_bitmap32[y_32][31-x_32];
                        font_in =  Hin_bitmap32[y_32][31-x_32];
                    end
                    [134:165] : begin                  
                        x_32 = x_pixel - (134);
                        font_out = Iout_bitmap32[y_32][31-x_32];
                        font_in =  Iin_bitmap32[y_32][31-x_32];
                    end
                    [168:199] : begin                  
                        x_32 = x_pixel - (168);
                        font_out = Gout_bitmap32[y_32][31-x_32];
                        font_in =  Gin_bitmap32[y_32][31-x_32];
                    end
                    [202:233] : begin                  
                        x_32 = x_pixel - (202);
                        font_out = Hout_bitmap32[y_32][31-x_32];
                        font_in =  Hin_bitmap32[y_32][31-x_32];
                    end
                    //space
                    [264:295] : begin                  
                        x_32 = x_pixel - (264);
                        font_out = Sout_bitmap32[y_32][31-x_32];
                        font_in =  Sin_bitmap32[y_32][31-x_32];
                    end
                    [298:329] : begin                  
                        x_32 = x_pixel - (298);
                        font_out = Cout_bitmap32[y_32][31-x_32];
                        font_in =  Cin_bitmap32[y_32][31-x_32];
                    end
                    [332:363] : begin                  
                        x_32 = x_pixel - (332);
                        font_out = Oout_bitmap32[y_32][31-x_32];
                        font_in =  Oin_bitmap32[y_32][31-x_32];
                    end
                    [366:397] : begin                  
                        x_32 = x_pixel - (366);
                        font_out = Rout_bitmap32[y_32][31-x_32];
                        font_in =  Rin_bitmap32[y_32][31-x_32];
                    end
                    [400:431] : begin                  
                        x_32 = x_pixel - (400);
                        font_out = Eout_bitmap32[y_32][31-x_32];
                        font_in =  Ein_bitmap32[y_32][31-x_32];
                    end
                    [434:465] : begin                  
                        x_32 = x_pixel - (434);
                        font_out = co_bitmapout_32[y_32][31-x_32];
                        font_in =  co_bitmapin_32[y_32][31-x_32];
                    end
                    [468:499] : begin   // high score          
                        x_32 = x_pixel - (468);
                        case (high_score / 10)
                        4'd0: begin
                            font_out = zeroout_bitmap32[y_32][31-x_32];
                            font_in = zeroin_bitmap32[y_32][31-x_32];
                        end 
                        4'd1: begin
                            font_out = oneout_bitmap32[y_32][31-x_32];
                            font_in = onein_bitmap32[y_32][31-x_32];
                        end 
                        4'd2: begin
                            font_out = twoout_bitmap32[y_32][31-x_32];
                            font_in = twoin_bitmap32[y_32][31-x_32];
                        end 
                        4'd3: begin
                            font_out = threeout_bitmap32[y_32][31-x_32];
                            font_in = threein_bitmap32[y_32][31-x_32];
                        end 
                        4'd4: begin
                            font_out = fourout_bitmap32[y_32][31-x_32];
                            font_in = fourin_bitmap32[y_32][31-x_32];
                        end 
                        4'd5: begin
                            font_out = fiveout_bitmap32[y_32][31-x_32];
                            font_in = fivein_bitmap32[y_32][31-x_32];
                        end 
                        4'd6: begin
                            font_out = sixout_bitmap32[y_32][31-x_32];
                            font_in = sixin_bitmap32[y_32][31-x_32];
                        end 
                        4'd7: begin
                            font_out = sevenout_bitmap32[y_32][31-x_32];
                            font_in = sevenin_bitmap32[y_32][31-x_32];
                        end 
                        4'd8: begin
                            font_out = eightout_bitmap32[y_32][31-x_32];
                            font_in = eightin_bitmap32[y_32][31-x_32];
                        end 
                        4'd9: begin
                            font_out = nineout_bitmap32[y_32][31-x_32];
                            font_in = ninein_bitmap32[y_32][31-x_32];
                        end 
                        endcase
                    end
                    [502:533] : begin   //high score               
                        x_32 = x_pixel - (502);
                        case (high_score % 10)
                        4'd0: begin
                            font_out = zeroout_bitmap32[y_32][31-x_32];
                            font_in = zeroin_bitmap32[y_32][31-x_32];
                        end 
                        4'd1: begin
                            font_out = oneout_bitmap32[y_32][31-x_32];
                            font_in = onein_bitmap32[y_32][31-x_32];
                        end 
                        4'd2: begin
                            font_out = twoout_bitmap32[y_32][31-x_32];
                            font_in = twoin_bitmap32[y_32][31-x_32];
                        end 
                        4'd3: begin
                            font_out = threeout_bitmap32[y_32][31-x_32];
                            font_in = threein_bitmap32[y_32][31-x_32];
                        end 
                        4'd4: begin
                            font_out = fourout_bitmap32[y_32][31-x_32];
                            font_in = fourin_bitmap32[y_32][31-x_32];
                        end 
                        4'd5: begin
                            font_out = fiveout_bitmap32[y_32][31-x_32];
                            font_in = fivein_bitmap32[y_32][31-x_32];
                        end 
                        4'd6: begin
                            font_out = sixout_bitmap32[y_32][31-x_32];
                            font_in = sixin_bitmap32[y_32][31-x_32];
                        end 
                        4'd7: begin
                            font_out = sevenout_bitmap32[y_32][31-x_32];
                            font_in = sevenin_bitmap32[y_32][31-x_32];
                        end 
                        4'd8: begin
                            font_out = eightout_bitmap32[y_32][31-x_32];
                            font_in = eightin_bitmap32[y_32][31-x_32];
                        end 
                        4'd9: begin
                            font_out = nineout_bitmap32[y_32][31-x_32];
                            font_in = ninein_bitmap32[y_32][31-x_32];
                        end 
                        endcase
                    end
                    endcase
                end else if (y_pixel >= 410 && y_pixel< 432) begin
                    y_32 = y_pixel - 410;
                    if (x_pixel >= 30 && x_pixel < 52) begin
                        x_32 = x_pixel - 30;
                        cha_1 = black[y_32][21-x_32];
                        cha_2 = white[y_32][21-x_32];
                        cha_3 = green[y_32][21-x_32];
                        cha_4 = lime[y_32][21-x_32];
                        cha_5 = skin[y_32][21-x_32];
                        cha_6 = pink[y_32][21-x_32];
                        cha_7 = yellow[y_32][21-x_32];
                    end
                end

                //sw = !q_start
                if (start_ff2) begin
                    state_next = START;
                end
            end


        START : begin 
                if (y_pixel >= RUNFORCOLOR_Y && y_pixel < RUNFORCOLOR_Y + SPACE_32 ) begin 
                    y_32 = y_pixel - RUNFORCOLOR_Y;

                    case (x_pixel) inside
                    [(RUNFORCOLOR_X):(RUNFORCOLOR_X + BIT31)] : begin //  100 ~ 131                  
                        x_32 = x_pixel - (RUNFORCOLOR_X);
                        font_out = Rout_bitmap32[y_32][31-x_32];
                        font_in = Rin_bitmap32[y_32][31-x_32];
                    end
                    [(RUNFORCOLOR_X + BIT31 + SPACE_3):(RUNFORCOLOR_X + 2*BIT31 + SPACE_3)] : begin //  134 ~ 165
                        x_32 = x_pixel - (RUNFORCOLOR_X+ BIT31 +SPACE_3);
                        font_out = Uout_bitmap32[y_32][31-x_32];
                        font_in = Uin_bitmap32[y_32][31-x_32];
                    end 
                    [(RUNFORCOLOR_X + 2*BIT31 + 2*SPACE_3):(RUNFORCOLOR_X + 3*BIT31 + 2*SPACE_3)] : begin // 168 ~ 199
                        x_32 = x_pixel - (RUNFORCOLOR_X + 2*BIT31 + 2*SPACE_3);
                        font_out = Nout_bitmap32[y_32][31-x_32];
                        font_in = Nin_bitmap32[y_32][31-x_32];
                    end
                    //space32
                    [(RUNFORCOLOR_X + 3*BIT31 + 3*SPACE_3 + SPACE_32):(RUNFORCOLOR_X + 4*BIT31 + 3*SPACE_3 + SPACE_32)] : begin // 168 ~ 199
                        x_32 = x_pixel - (RUNFORCOLOR_X + 3*BIT31 + 3*SPACE_3 + SPACE_32);
                        font_out = Fout_bitmap32[y_32][31-x_32];
                        font_in = Fin_bitmap32[y_32][31-x_32];
                    end
                    [(RUNFORCOLOR_X + 4*BIT31 + 4*SPACE_3 + SPACE_32):(RUNFORCOLOR_X + 5*BIT31 + 4*SPACE_3 + SPACE_32)] : begin // 168 ~ 199
                        x_32 = x_pixel - (RUNFORCOLOR_X + 4*BIT31 + 4*SPACE_3 + SPACE_32);
                        font_out = Oout_bitmap32[y_32][31-x_32];
                        font_in = Oin_bitmap32[y_32][31-x_32];
                    end
                    [(RUNFORCOLOR_X + 5*BIT31 + 5*SPACE_3 + SPACE_32):(RUNFORCOLOR_X + 6*BIT31 + 5*SPACE_3 + SPACE_32)] : begin // 168 ~ 199
                        x_32 = x_pixel - (RUNFORCOLOR_X + 5*BIT31 + 5*SPACE_3 + SPACE_32);
                        font_out = Rout_bitmap32[y_32][31-x_32];
                        font_in = Rin_bitmap32[y_32][31-x_32];
                    end
                    //space32
                    [(RUNFORCOLOR_X + 6*BIT31 + 6*SPACE_3 + 2*SPACE_32):(RUNFORCOLOR_X + 7*BIT31 + 6*SPACE_3 + 2*SPACE_32)] : begin // 168 ~ 199
                        x_32 = x_pixel - (RUNFORCOLOR_X + 6*BIT31 + 6*SPACE_3 + 2*SPACE_32);
                        font_out = Cout_bitmap32[y_32][31-x_32];
                        font_in = Cin_bitmap32[y_32][31-x_32];
                    end
                    [(RUNFORCOLOR_X + 7*BIT31 + 7*SPACE_3 + 2*SPACE_32):(RUNFORCOLOR_X + 8*BIT31 + 7*SPACE_3 + 2*SPACE_32)] : begin // 168 ~ 199
                        x_32 = x_pixel - (RUNFORCOLOR_X + 7*BIT31 + 7*SPACE_3 + 2*SPACE_32);
                        font_out = Oout_bitmap32[y_32][31-x_32];
                        font_in = Oin_bitmap32[y_32][31-x_32];
                    end
                    [(RUNFORCOLOR_X + 8*BIT31 + 8*SPACE_3 + 2*SPACE_32):(RUNFORCOLOR_X + 9*BIT31 + 8*SPACE_3 + 2*SPACE_32)] : begin // 168 ~ 199
                        x_32 = x_pixel - (RUNFORCOLOR_X + 8*BIT31 + 8*SPACE_3 + 2*SPACE_32);
                        font_out = Lout_bitmap32[y_32][31-x_32];
                        font_in = Lin_bitmap32[y_32][31-x_32];
                    end
                    [(RUNFORCOLOR_X + 9*BIT31 + 9*SPACE_3 + 2*SPACE_32):(RUNFORCOLOR_X + 10*BIT31 + 9*SPACE_3 + 2*SPACE_32)] : begin // 168 ~ 199
                        x_32 = x_pixel - (RUNFORCOLOR_X + 9*BIT31 + 9*SPACE_3 + 2*SPACE_32);
                        font_out = Oout_bitmap32[y_32][31-x_32];
                        font_in = Oin_bitmap32[y_32][31-x_32];
                    end
                    [(RUNFORCOLOR_X + 10*BIT31 + 10*SPACE_3 + 2*SPACE_32):(RUNFORCOLOR_X + 11*BIT31 + 10*SPACE_3 + 2*SPACE_32)] : begin // 168 ~ 199
                        x_32 = x_pixel - (RUNFORCOLOR_X + 10*BIT31 + 10*SPACE_3 + 2*SPACE_32);
                        font_out = Rout_bitmap32[y_32][31-x_32];
                        font_in = Rin_bitmap32[y_32][31-x_32];
                    end
                    endcase
                end    

                // 3,2,1,0 표시
                else if (y_pixel >= 136 && y_pixel < 136 + SPACE_32) begin
                    y_32 = y_pixel - 136;
                    if (x_pixel >= 420 && x_pixel < 420 + SPACE_32) begin
                        x_32 = x_pixel - 420;
                        case (startcount)
                            2'd0: begin
                                font_out = zeroout_bitmap32[y_32][31-x_32];
                                font_in  = zeroin_bitmap32[y_32][31-x_32];
                            end 
                            2'd1: begin
                                font_out = oneout_bitmap32[y_32][31-x_32];
                                font_in  = onein_bitmap32[y_32][31-x_32];
                            end 
                            2'd2: begin
                                font_out = twoout_bitmap32[y_32][31-x_32];
                                font_in  = twoin_bitmap32[y_32][31-x_32];
                            end 
                            2'd3: begin
                                font_out = threeout_bitmap32[y_32][31-x_32];
                                font_in  = threein_bitmap32[y_32][31-x_32];
                            end 
                        endcase
                    end
                end


            if (clk_counter == 25_000_000 - 1) begin
                clk_counter_next = 0;  // 카운터 초기화
                if (startcount > 0) begin
                    startcount_next = startcount - 1;  // 카운트다운 감소
                end else begin
                    startcount_next = 0;  // 카운트다운이 0이 되면 유지
                    state_next = LEVEL0;
                end
            end else begin
                clk_counter_next = clk_counter + 1;  // 카운터 증가
            end
        end

        /************************************LEVEL0******************************************/
        /************************************LEVEL0******************************************/
        /************************************LEVEL0******************************************/
        /************************************LEVEL0******************************************/
        /************************************LEVEL0******************************************/
        /************************************LEVEL0******************************************/
        /************************************LEVEL0******************************************/
        /************************************LEVEL0******************************************/
        /************************************LEVEL0******************************************/
        /************************************LEVEL0******************************************/



            LEVEL0: // 연습 게임, 색깔 1개 보여주고, win/lose 판별
            begin
                // 문제에 따라 색깔 1개 표시, (y= 80~200, x= 260 ~ 380) 
                lvl_count_next = 0;     // 레벨 카운터 초기화
                game_done_next = 1;
                led_next = 4'b0001;
                if ((x_pixel < 380 && x_pixel >= 260) && (y_pixel < 200 && y_pixel >= 80)) begin
                    case (question[1:0])
                        2'd0: {red_port, green_port, blue_port} = {4'h0, 4'h0, 4'h0}; //black, 0 들어오면 검정색
                        2'd1: {red_port, green_port, blue_port} = {4'hf, 4'h0, 4'h0}; //red
                        2'd2: {red_port, green_port, blue_port} = {4'hf, 4'hf, 4'h0}; //yellow
                        2'd3: {red_port, green_port, blue_port} = {4'h0, 4'h0, 4'hf}; //blue
                    endcase   
                end
                // 정답 맞힐 수 있는 영역 표시(검정색)    (y= 280~400, x= 260 ~ 380)   
                else if (((x_pixel < 380 && x_pixel >= 260) && (y_pixel == 280 || y_pixel == 400)) ||
                        ((x_pixel == 380 || x_pixel == 260) && (y_pixel >= 280 && y_pixel < 400))) begin
                        red_port   = 4'h0;  // Red
                        green_port = 4'h0;  // Green
                        blue_port  = 4'h0;  // Blue  
                end


                // LEVEL 0 표시     (y= 28~60, x= 210 ~ 436)
                else if (y_pixel >= 28 && y_pixel < 60) begin
                    y_32 = y_pixel - 28;
                    case (x_pixel) inside
                        [210:241]: begin        // L
                            x_32 = x_pixel - (210);
                            font_out = Lout_bitmap32[y_32][31-x_32];
                            font_in = Lin_bitmap32[y_32][31-x_32];
                        end
                        [243:274]: begin        // E
                            x_32 = x_pixel - (243);
                            font_out = Eout_bitmap32[y_32][31-x_32];
                            font_in = Ein_bitmap32[y_32][31-x_32];
                        end
                        [276:307]: begin        // V
                            x_32 = x_pixel - (276);
                            font_out = Vout_bitmap32[y_32][31-x_32];
                            font_in = Vin_bitmap32[y_32][31-x_32];
                        end
                        [309:340]: begin        // E
                            x_32 = x_pixel - (309);
                            font_out = Eout_bitmap32[y_32][31-x_32];
                            font_in = Ein_bitmap32[y_32][31-x_32];
                        end
                        [342:373]: begin        // L
                            x_32 = x_pixel - (342);
                            font_out = Lout_bitmap32[y_32][31-x_32];
                            font_in = Lin_bitmap32[y_32][31-x_32];
                        end
                        [405:436]: begin        // 0
                            x_32 = x_pixel - (405);
                            font_out = zeroout_bitmap32[y_32][31-x_32];
                            font_in = zeroin_bitmap32[y_32][31-x_32];
                        end
                        [550:581]: begin       // countdown (y= 28~60, x=500~532 )
                            x_32 = x_pixel - (550);
                            case (countdown)
                            4'd0: begin
                                font_out = zeroout_bitmap32[y_32][31-x_32];
                                countcolor_in = zeroin_bitmap32[y_32][31-x_32];
                            end 
                            4'd1: begin
                                font_out = oneout_bitmap32[y_32][31-x_32];
                                countcolor_in = onein_bitmap32[y_32][31-x_32];
                            end 
                            4'd2: begin
                                font_out = twoout_bitmap32[y_32][31-x_32];
                                countcolor_in = twoin_bitmap32[y_32][31-x_32];
                            end 
                            4'd3: begin
                                font_out = threeout_bitmap32[y_32][31-x_32];
                                countcolor_in = threein_bitmap32[y_32][31-x_32];
                            end 
                            4'd4: begin
                                font_out = fourout_bitmap32[y_32][31-x_32];
                                countcolor_in = fourin_bitmap32[y_32][31-x_32];
                            end 
                            4'd5: begin
                                font_out = fiveout_bitmap32[y_32][31-x_32];
                                countcolor_in = fivein_bitmap32[y_32][31-x_32];
                            end 
                            4'd6: begin
                                font_out = sixout_bitmap32[y_32][31-x_32];
                                countcolor_in = sixin_bitmap32[y_32][31-x_32];
                            end 
                            4'd7: begin
                                font_out = sevenout_bitmap32[y_32][31-x_32];
                                countcolor_in = sevenin_bitmap32[y_32][31-x_32];
                            end 
                            4'd8: begin
                                font_out = eightout_bitmap32[y_32][31-x_32];
                                countcolor_in = eightin_bitmap32[y_32][31-x_32];
                            end 
                            4'd9: begin
                                font_out = nineout_bitmap32[y_32][31-x_32];
                                countcolor_in = ninein_bitmap32[y_32][31-x_32];
                            end 
                            endcase
                        end
                    endcase
                end

          



                // 카운트다운을 위한 카운터
                if (clk_counter == 25_000_000 - 1) begin
                    clk_counter_next = 0;  // 카운터 초기화
                    if (countdown > 0) begin
                        countdown_next = countdown - 1;  // 카운트다운 감소
                    end else begin
                        countdown_next = 0;  // 카운트다운이 0이 되면 유지
                    end
                end else begin
                    clk_counter_next = clk_counter + 1;  // 카운터 증가
                end






                // 카운트다운 후에 win/lose 디스플레이 표시
                if (countdown == 0) begin
                    //win_lose가 안들어오면 계속 1을 주는 문제 발생?
                    countdown_done_next = 1;  // 카운트다운 완료 신호
                    state_next = WIN_LOSE;
                end 
            end




        /************************************LEVEL1-1******************************************/
        /************************************LEVEL1-1******************************************/
        /************************************LEVEL1-1******************************************/
        /************************************LEVEL1-1******************************************/
        /************************************LEVEL1-1******************************************/
        /************************************LEVEL1-1******************************************/
        /************************************LEVEL1-1******************************************/
        /************************************LEVEL1-1******************************************/
        /************************************LEVEL1-1******************************************/
        /************************************LEVEL1-1******************************************/
            LEVEL1_1: // 깜빡 + 색 2개 표시 
            begin
                game_done_next = 1;
                // 0.2초 마다 깜빡 
                led_next = 4'b0010;
                if (clk_counter_blink == 5_000_000 - 1) begin
                    clk_counter_blink_next = 0;  // 카운터 초기화
                    if (blink_count == 49) begin
                        blink_count_next = 0;
                    end else begin
                        blink_count_next = blink_count + 1;
                    end

                end else begin
                    clk_counter_blink_next = clk_counter_blink + 1;  // 카운터 증가
                end



                // 0.2~0.4초 처음 색 보여줌, 0.6~0.8초 두번째 색 보여줌, (y= 80~200, x= 260 ~ 380) 
                if ((x_pixel < 380 && x_pixel >= 260) && (y_pixel < 200 && y_pixel >= 80)) begin      
                    case (blink_count)
                        6'd1: begin
                            case (question[1:0])
                            2'd0: {red_port, green_port, blue_port} = {4'h0, 4'h0, 4'h0}; //black, 0 들어오면 검정색
                            2'd1: {red_port, green_port, blue_port} = {4'hf, 4'h0, 4'h0}; //red
                            2'd2: {red_port, green_port, blue_port} = {4'hf, 4'hf, 4'h0}; //yellow
                            2'd3: {red_port, green_port, blue_port} = {4'h0, 4'h0, 4'hf}; //blue
                        endcase
                        end
                        6'd3: begin
                            q_display_done_next = 1;
                            case (question[3:2])
                            2'd0: {red_port, green_port, blue_port} = {4'h0, 4'h0, 4'h0}; //black
                            2'd1: {red_port, green_port, blue_port} = {4'hf, 4'h0, 4'h0}; //red
                            2'd2: {red_port, green_port, blue_port} = {4'hf, 4'hf, 4'h0}; //yellow
                            2'd3: {red_port, green_port, blue_port} = {4'h0, 4'h0, 4'hf}; //blue
                        endcase
                        end
                        default: begin
                            {red_port, green_port, blue_port} = {cam_r, cam_g, cam_b}; // 깜빡이지 않을떈 아무것도 표시 X
                        end
                    endcase
                end  
                   

                 // 정답 제출할 영역 표시 (검정색) , (y= 280~400, x= 150 ~ 270), (y= 280~400, x= 370 ~ 490)  
                else if (((x_pixel < 270 && x_pixel >= 150) && (y_pixel == 280 || y_pixel == 400)) ||
                        ((x_pixel == 270 || x_pixel == 150) && (y_pixel >= 280 && y_pixel < 400))) begin
                    red_port   = 4'h0;  // Red
                    green_port = 4'h0;  // Green
                    blue_port  = 4'h0;  // Blue  
                end else if (((x_pixel < 490 && x_pixel >= 370) && (y_pixel == 280 || y_pixel == 400)) ||
                        ((x_pixel == 490 || x_pixel == 370) && (y_pixel >= 280 && y_pixel < 400))) begin
                    red_port   = 4'h0;  // Red
                    green_port = 4'h0;  // Green
                    blue_port  = 4'h0;  // Blue  
                end

                // LEVEL 1-1 표시     (y= 28~60, x= 210 ~ 436) 
                else if (y_pixel >= 28 && y_pixel < 60) begin
                    y_32 = y_pixel - 28;
                    case (x_pixel) inside
                        [210:241]: begin        // L
                            x_32 = x_pixel - (210);
                            font_out = Lout_bitmap32[y_32][31-x_32];
                            font_in = Lin_bitmap32[y_32][31-x_32];
                        end
                        [243:274]: begin        // E
                            x_32 = x_pixel - (243);
                            font_out = Eout_bitmap32[y_32][31-x_32];
                            font_in = Ein_bitmap32[y_32][31-x_32];
                        end
                        [276:307]: begin        // V
                            x_32 = x_pixel - (276);
                            font_out = Vout_bitmap32[y_32][31-x_32];
                            font_in = Vin_bitmap32[y_32][31-x_32];
                        end
                        [309:340]: begin        // E
                            x_32 = x_pixel - (309);
                            font_out = Eout_bitmap32[y_32][31-x_32];
                            font_in = Ein_bitmap32[y_32][31-x_32];
                        end
                        [342:373]: begin        // L
                            x_32 = x_pixel - (342);
                            font_out = Lout_bitmap32[y_32][31-x_32];
                            font_in = Lin_bitmap32[y_32][31-x_32];
                        end
                        [405:436]: begin        // 1
                            x_32 = x_pixel - (405);
                            font_out = oneout_bitmap32[y_32][31-x_32];
                            font_in = onein_bitmap32[y_32][31-x_32];
                        end
                        [440:471]: begin        // -
                            x_32 = x_pixel - (440);
                            font_out = dashout_bitmap32[y_32][31-x_32];
                            font_in = dashin_bitmap32[y_32][31-x_32];
                        end
                        [475:506]: begin        // 1
                            x_32 = x_pixel - (475);
                            font_out = oneout_bitmap32[y_32][31-x_32];
                            font_in = onein_bitmap32[y_32][31-x_32];
                        end
                        [550:581]: begin       // countdown (y= 28~60, x=500~532 )
                        if (q_display_done) begin
                            x_32 = x_pixel - (550);
                            case (countdown)
                            4'd0: begin
                                font_out = zeroout_bitmap32[y_32][31-x_32];
                                countcolor_in = zeroin_bitmap32[y_32][31-x_32];
                            end 
                            4'd1: begin
                                font_out = oneout_bitmap32[y_32][31-x_32];
                                countcolor_in = onein_bitmap32[y_32][31-x_32];
                            end 
                            4'd2: begin
                                font_out = twoout_bitmap32[y_32][31-x_32];
                                countcolor_in = twoin_bitmap32[y_32][31-x_32];
                            end 
                            4'd3: begin
                                font_out = threeout_bitmap32[y_32][31-x_32];
                                countcolor_in = threein_bitmap32[y_32][31-x_32];
                            end 
                            4'd4: begin
                                font_out = fourout_bitmap32[y_32][31-x_32];
                                countcolor_in = fourin_bitmap32[y_32][31-x_32];
                            end 
                            4'd5: begin
                                font_out = fiveout_bitmap32[y_32][31-x_32];
                                countcolor_in = fivein_bitmap32[y_32][31-x_32];
                            end 
                            4'd6: begin
                                font_out = sixout_bitmap32[y_32][31-x_32];
                                countcolor_in = sixin_bitmap32[y_32][31-x_32];
                            end 
                            4'd7: begin
                                font_out = sevenout_bitmap32[y_32][31-x_32];
                                countcolor_in = sevenin_bitmap32[y_32][31-x_32];
                            end 
                            4'd8: begin
                                font_out = eightout_bitmap32[y_32][31-x_32];
                                countcolor_in = eightin_bitmap32[y_32][31-x_32];
                            end 
                            4'd9: begin
                                font_out = nineout_bitmap32[y_32][31-x_32];
                                countcolor_in = ninein_bitmap32[y_32][31-x_32];
                            end 
                            endcase
                        end
                        end
                    endcase
                end


                // 카운트다운용 카운터 
                if (clk_counter == 25_000_000 - 1) begin
                    clk_counter_next = 0;  // 카운터 초기화
                    if (countdown > 0) begin
                        countdown_next = countdown - 1;  // 카운트다운 감소
                    end else begin
                        countdown_next = 0;  // 카운트다운이 0이 되면 유지
                    end
                end else begin
                    clk_counter_next = clk_counter + 1;  // 카운터 증가
                end


                if (countdown == 0) begin
                    countdown_done_next = 1;  // 카운트다운 완료 신호
                    q_display_done_next = 0;
                    state_next = WIN_LOSE;        
                end 
            end

        /************************************LEVEL1-2******************************************/
        /************************************LEVEL1-2******************************************/
        /************************************LEVEL1-2******************************************/
        /************************************LEVEL1-2******************************************/
        /************************************LEVEL1-2******************************************/
        /************************************LEVEL1-2******************************************/
        /************************************LEVEL1-2******************************************/
        /************************************LEVEL1-2******************************************/
        /************************************LEVEL1-2******************************************/
        /************************************LEVEL1-2******************************************/
         LEVEL1_2: // 깜빡 + 색 3개 표시 
            begin
                game_done_next = 1;
                // 0.2초 마다 깜빡 
                led_next = 4'b0010;
                if (clk_counter_blink == 5_000_000 - 1) begin
                    clk_counter_blink_next = 0;  // 카운터 초기화
                    if (blink_count == 49) begin
                        blink_count_next = 0;
                    end else begin
                        blink_count_next = blink_count + 1;
                    end

                end else begin
                    clk_counter_blink_next = clk_counter_blink + 1;  // 카운터 증가
                end



                // 0.2~0.4초 처음 색 보여줌, 0.6~0.8초 두번째 색 보여줌, 1~1.2초 세번째 색 보여줌줌 (y= 80~200, x= 260 ~ 380) 
                if ((x_pixel < 380 && x_pixel >= 260) && (y_pixel < 200 && y_pixel >= 80)) begin      
                    case (blink_count)
                        6'd1: begin
                            case (question[1:0])
                            2'd0: {red_port, green_port, blue_port} = {4'h0, 4'h0, 4'h0}; //black, 0 들어오면 검정색
                            2'd1: {red_port, green_port, blue_port} = {4'hf, 4'h0, 4'h0}; //red
                            2'd2: {red_port, green_port, blue_port} = {4'hf, 4'hf, 4'h0}; //yellow
                            2'd3: {red_port, green_port, blue_port} = {4'h0, 4'h0, 4'hf}; //blue
                        endcase
                        end
                        6'd3: begin
                            case (question[3:2])
                            2'd0: {red_port, green_port, blue_port} = {4'h0, 4'h0, 4'h0}; //black
                            2'd1: {red_port, green_port, blue_port} = {4'hf, 4'h0, 4'h0}; //red
                            2'd2: {red_port, green_port, blue_port} = {4'hf, 4'hf, 4'h0}; //yellow
                            2'd3: {red_port, green_port, blue_port} = {4'h0, 4'h0, 4'hf}; //blue
                        endcase
                        end
                        6'd5: begin
                            q_display_done_next = 1;
                            case (question[5:4])
                            2'd0: {red_port, green_port, blue_port} = {4'h0, 4'h0, 4'h0}; //black
                            2'd1: {red_port, green_port, blue_port} = {4'hf, 4'h0, 4'h0}; //red
                            2'd2: {red_port, green_port, blue_port} = {4'hf, 4'hf, 4'h0}; //yellow
                            2'd3: {red_port, green_port, blue_port} = {4'h0, 4'h0, 4'hf}; //blue
                        endcase
                        end
                        default: begin
                            {red_port, green_port, blue_port} = {cam_r, cam_g, cam_b}; // 깜빡이지 않을떈 아무것도 표시 X
                        end
                    endcase
                end  
                   

                // 정답 제출할 영역 표시 (y= 280~400, x= 70 ~ 190), (y= 280~400, x= 260 ~ 380) , (y= 280~400, x= 450 ~ 570)  
                else if (((x_pixel < 190 && x_pixel >= 70) && (y_pixel == 280 || y_pixel == 400)) ||
                        ((x_pixel == 190 || x_pixel == 70) && (y_pixel >= 280 && y_pixel < 400))) begin
                    red_port   = 4'h0;  
                    green_port = 4'h0;  
                    blue_port  = 4'h0;  // -> black 
                end else if (((x_pixel < 380 && x_pixel >= 260) && (y_pixel == 280 || y_pixel == 400)) ||
                        ((x_pixel == 380 || x_pixel == 260) && (y_pixel >= 280 && y_pixel < 400))) begin
                    red_port   = 4'h0;  
                    green_port = 4'h0;  
                    blue_port  = 4'h0;  // -> black  
                end else if (((x_pixel < 570 && x_pixel >= 450) && (y_pixel == 280 || y_pixel == 400)) ||
                        ((x_pixel == 570 || x_pixel == 450) && (y_pixel >= 280 && y_pixel < 400))) begin
                    red_port   = 4'h0;  
                    green_port = 4'h0;  
                    blue_port  = 4'h0;  // -> black  
                end 

                // LEVEL 1-2 표시     (y= 28~60, x= 210 ~ 436) 
                else if (y_pixel >= 28 && y_pixel < 60) begin
                    y_32 = y_pixel - 28;
                    case (x_pixel) inside
                        [210:241]: begin        // L
                            x_32 = x_pixel - (210);
                            font_out = Lout_bitmap32[y_32][31-x_32];
                            font_in = Lin_bitmap32[y_32][31-x_32];
                        end
                        [243:274]: begin        // E
                            x_32 = x_pixel - (243);
                            font_out = Eout_bitmap32[y_32][31-x_32];
                            font_in = Ein_bitmap32[y_32][31-x_32];
                        end
                        [276:307]: begin        // V
                            x_32 = x_pixel - (276);
                            font_out = Vout_bitmap32[y_32][31-x_32];
                            font_in = Vin_bitmap32[y_32][31-x_32];
                        end
                        [309:340]: begin        // E
                            x_32 = x_pixel - (309);
                            font_out = Eout_bitmap32[y_32][31-x_32];
                            font_in = Ein_bitmap32[y_32][31-x_32];
                        end
                        [342:373]: begin        // L
                            x_32 = x_pixel - (342);
                            font_out = Lout_bitmap32[y_32][31-x_32];
                            font_in = Lin_bitmap32[y_32][31-x_32];
                        end
                        [405:436]: begin        // 1
                            x_32 = x_pixel - (405);
                            font_out = oneout_bitmap32[y_32][31-x_32];
                            font_in = onein_bitmap32[y_32][31-x_32];
                        end
                        [440:471]: begin        // -
                            x_32 = x_pixel - (440);
                            font_out = dashout_bitmap32[y_32][31-x_32];
                            font_in = dashin_bitmap32[y_32][31-x_32];
                        end
                        [475:506]: begin        // 2
                            x_32 = x_pixel - (475);
                            font_out = twoout_bitmap32[y_32][31-x_32];
                            font_in = twoin_bitmap32[y_32][31-x_32];
                        end
                        [550:581]: begin       // countdown (y= 28~60, x=500~532 )
                        if (q_display_done) begin
                            x_32 = x_pixel - (550);
                            case (countdown)
                            4'd0: begin
                                font_out = zeroout_bitmap32[y_32][31-x_32];
                                countcolor_in = zeroin_bitmap32[y_32][31-x_32];
                            end 
                            4'd1: begin
                                font_out = oneout_bitmap32[y_32][31-x_32];
                                countcolor_in = onein_bitmap32[y_32][31-x_32];
                            end 
                            4'd2: begin
                                font_out = twoout_bitmap32[y_32][31-x_32];
                                countcolor_in = twoin_bitmap32[y_32][31-x_32];
                            end 
                            4'd3: begin
                                font_out = threeout_bitmap32[y_32][31-x_32];
                                countcolor_in = threein_bitmap32[y_32][31-x_32];
                            end 
                            4'd4: begin
                                font_out = fourout_bitmap32[y_32][31-x_32];
                                countcolor_in = fourin_bitmap32[y_32][31-x_32];
                            end 
                            4'd5: begin
                                font_out = fiveout_bitmap32[y_32][31-x_32];
                                countcolor_in = fivein_bitmap32[y_32][31-x_32];
                            end 
                            4'd6: begin
                                font_out = sixout_bitmap32[y_32][31-x_32];
                                countcolor_in = sixin_bitmap32[y_32][31-x_32];
                            end 
                            4'd7: begin
                                font_out = sevenout_bitmap32[y_32][31-x_32];
                                countcolor_in = sevenin_bitmap32[y_32][31-x_32];
                            end 
                            4'd8: begin
                                font_out = eightout_bitmap32[y_32][31-x_32];
                                countcolor_in = eightin_bitmap32[y_32][31-x_32];
                            end 
                            4'd9: begin
                                font_out = nineout_bitmap32[y_32][31-x_32];
                                countcolor_in = ninein_bitmap32[y_32][31-x_32];
                            end 
                            endcase
                        end
                        end
                    endcase
                end


                // 카운트다운용 카운터 
                if (clk_counter == 25_000_000 - 1) begin
                    clk_counter_next = 0;  // 카운터 초기화
                    if (countdown > 0) begin
                        countdown_next = countdown - 1;  // 카운트다운 감소
                    end else begin
                        countdown_next = 0;  // 카운트다운이 0이 되면 유지
                    end
                end else begin
                    clk_counter_next = clk_counter + 1;  // 카운터 증가
                end


                if (countdown == 0) begin
                    countdown_done_next = 1;  // 카운트다운 완료 신호
                    q_display_done_next = 0;
                    state_next = WIN_LOSE;        
                end 
            end


        

        /************************************LEVEL1-3******************************************/
        /************************************LEVEL1-3******************************************/
        /************************************LEVEL1-3******************************************/
        /************************************LEVEL1-3******************************************/
        /************************************LEVEL1-3******************************************/
        /************************************LEVEL1-3******************************************/
        /************************************LEVEL1-3******************************************/
        /************************************LEVEL1-3******************************************/
        /************************************LEVEL1-3******************************************/
        /************************************LEVEL1-3******************************************/
         LEVEL1_3: // 깜빡 + 색 4개 표시 
            begin
                game_done_next = 1;
                // 0.2초 마다 깜빡 
                led_next = 4'b0010;
                if (clk_counter_blink == 5_000_000 - 1) begin
                    clk_counter_blink_next = 0;  // 카운터 초기화
                    if (blink_count == 49) begin
                        blink_count_next = 0;
                    end else begin
                        blink_count_next = blink_count + 1;
                    end

                end else begin
                    clk_counter_blink_next = clk_counter_blink + 1;  // 카운터 증가
                end



                // 0.2~0.4초 처음 색 보여줌, 0.6~0.8초 두번째 색 보여줌, (y= 80~200, x= 260 ~ 380) 
                if ((x_pixel < 380 && x_pixel >= 260) && (y_pixel < 200 && y_pixel >= 80)) begin      
                    case (blink_count)
                        6'd1: begin
                            case (question[1:0])
                            2'd0: {red_port, green_port, blue_port} = {4'h0, 4'h0, 4'h0}; //black, 0 들어오면 검정색
                            2'd1: {red_port, green_port, blue_port} = {4'hf, 4'h0, 4'h0}; //red
                            2'd2: {red_port, green_port, blue_port} = {4'hf, 4'hf, 4'h0}; //yellow
                            2'd3: {red_port, green_port, blue_port} = {4'h0, 4'h0, 4'hf}; //blue
                        endcase
                        end
                        6'd3: begin
                            case (question[3:2])
                            2'd0: {red_port, green_port, blue_port} = {4'h0, 4'h0, 4'h0}; //black
                            2'd1: {red_port, green_port, blue_port} = {4'hf, 4'h0, 4'h0}; //red
                            2'd2: {red_port, green_port, blue_port} = {4'hf, 4'hf, 4'h0}; //yellow
                            2'd3: {red_port, green_port, blue_port} = {4'h0, 4'h0, 4'hf}; //blue
                        endcase
                        end
                        6'd5: begin
                            case (question[5:4])
                            2'd0: {red_port, green_port, blue_port} = {4'h0, 4'h0, 4'h0}; //black
                            2'd1: {red_port, green_port, blue_port} = {4'hf, 4'h0, 4'h0}; //red
                            2'd2: {red_port, green_port, blue_port} = {4'hf, 4'hf, 4'h0}; //yellow
                            2'd3: {red_port, green_port, blue_port} = {4'h0, 4'h0, 4'hf}; //blue
                        endcase
                        end
                        6'd7: begin
                            q_display_done_next = 1;
                            case (question[7:6])
                            2'd0: {red_port, green_port, blue_port} = {4'h0, 4'h0, 4'h0}; //black
                            2'd1: {red_port, green_port, blue_port} = {4'hf, 4'h0, 4'h0}; //red
                            2'd2: {red_port, green_port, blue_port} = {4'hf, 4'hf, 4'h0}; //yellow
                            2'd3: {red_port, green_port, blue_port} = {4'h0, 4'h0, 4'hf}; //blue
                        endcase
                        end
                        default: begin
                            {red_port, green_port, blue_port} = {cam_r, cam_g, cam_b}; // 깜빡이지 않을떈 아무것도 표시 X
                        end
                    endcase
                end  
                   

                // 정답 제출할 영역 표시 (y= 280~400, x= 32 ~ 152), (y= 280~400, x= 184 ~ 304) , (y= 280~400, x= 336 ~ 456)  , (y= 280~400, x= 488 ~ 608)  
                else if (((x_pixel < 152 && x_pixel >= 32) && (y_pixel == 280 || y_pixel == 400)) ||
                        ((x_pixel == 152 || x_pixel == 32) && (y_pixel >= 280 && y_pixel < 400))) begin
                    red_port   = 4'h0;  
                    green_port = 4'h0;  
                    blue_port  = 4'h0;  // -> black 
                end else if (((x_pixel < 304 && x_pixel >= 184) && (y_pixel == 280 || y_pixel == 400)) ||
                            ((x_pixel == 304 || x_pixel == 184) && (y_pixel >= 280 && y_pixel < 400))) begin
                    red_port   = 4'h0;  
                    green_port = 4'h0;  
                    blue_port  = 4'h0;  // -> black  
                end else if (((x_pixel < 456 && x_pixel >= 336) && (y_pixel == 280 || y_pixel == 400)) ||
                            ((x_pixel == 456 || x_pixel == 336) && (y_pixel >= 280 && y_pixel < 400))) begin
                    red_port   = 4'h0;  
                    green_port = 4'h0;  
                    blue_port  = 4'h0;  // -> black  
                end else if (((x_pixel < 608 && x_pixel >= 488) && (y_pixel == 280 || y_pixel == 400)) ||
                            ((x_pixel == 608 || x_pixel == 488) && (y_pixel >= 280 && y_pixel < 400))) begin
                    red_port   = 4'h0;  
                    green_port = 4'h0;  
                    blue_port  = 4'h0;  // -> black  
                end 


                // LEVEL 1-3 표시     (y= 28~60, x= 210 ~ 436) 
                else if (y_pixel >= 28 && y_pixel < 60) begin
                    y_32 = y_pixel - 28;
                    case (x_pixel) inside
                        [210:241]: begin        // L
                            x_32 = x_pixel - (210);
                            font_out = Lout_bitmap32[y_32][31-x_32];
                            font_in = Lin_bitmap32[y_32][31-x_32];
                        end
                        [243:274]: begin        // E
                            x_32 = x_pixel - (243);
                            font_out = Eout_bitmap32[y_32][31-x_32];
                            font_in = Ein_bitmap32[y_32][31-x_32];
                        end
                        [276:307]: begin        // V
                            x_32 = x_pixel - (276);
                            font_out = Vout_bitmap32[y_32][31-x_32];
                            font_in = Vin_bitmap32[y_32][31-x_32];
                        end
                        [309:340]: begin        // E
                            x_32 = x_pixel - (309);
                            font_out = Eout_bitmap32[y_32][31-x_32];
                            font_in = Ein_bitmap32[y_32][31-x_32];
                        end
                        [342:373]: begin        // L
                            x_32 = x_pixel - (342);
                            font_out = Lout_bitmap32[y_32][31-x_32];
                            font_in = Lin_bitmap32[y_32][31-x_32];
                        end
                        [405:436]: begin        // 1
                            x_32 = x_pixel - (405);
                            font_out = oneout_bitmap32[y_32][31-x_32];
                            font_in = onein_bitmap32[y_32][31-x_32];
                        end
                        [440:471]: begin        // -
                            x_32 = x_pixel - (440);
                            font_out = dashout_bitmap32[y_32][31-x_32];
                            font_in = dashin_bitmap32[y_32][31-x_32];
                        end
                        [475:506]: begin        // 3
                            x_32 = x_pixel - (475);
                            font_out = threeout_bitmap32[y_32][31-x_32];
                            font_in = threein_bitmap32[y_32][31-x_32];
                        end
                        [550:581]: begin       // countdown (y= 28~60, x=500~532 )
                        if (q_display_done) begin
                            x_32 = x_pixel - (550);
                            case (countdown)
                            4'd0: begin
                                font_out = zeroout_bitmap32[y_32][31-x_32];
                                countcolor_in = zeroin_bitmap32[y_32][31-x_32];
                            end 
                            4'd1: begin
                                font_out = oneout_bitmap32[y_32][31-x_32];
                                countcolor_in = onein_bitmap32[y_32][31-x_32];
                            end 
                            4'd2: begin
                                font_out = twoout_bitmap32[y_32][31-x_32];
                                countcolor_in = twoin_bitmap32[y_32][31-x_32];
                            end 
                            4'd3: begin
                                font_out = threeout_bitmap32[y_32][31-x_32];
                                countcolor_in = threein_bitmap32[y_32][31-x_32];
                            end 
                            4'd4: begin
                                font_out = fourout_bitmap32[y_32][31-x_32];
                                countcolor_in = fourin_bitmap32[y_32][31-x_32];
                            end 
                            4'd5: begin
                                font_out = fiveout_bitmap32[y_32][31-x_32];
                                countcolor_in = fivein_bitmap32[y_32][31-x_32];
                            end 
                            4'd6: begin
                                font_out = sixout_bitmap32[y_32][31-x_32];
                                countcolor_in = sixin_bitmap32[y_32][31-x_32];
                            end 
                            4'd7: begin
                                font_out = sevenout_bitmap32[y_32][31-x_32];
                                countcolor_in = sevenin_bitmap32[y_32][31-x_32];
                            end 
                            4'd8: begin
                                font_out = eightout_bitmap32[y_32][31-x_32];
                                countcolor_in = eightin_bitmap32[y_32][31-x_32];
                            end 
                            4'd9: begin
                                font_out = nineout_bitmap32[y_32][31-x_32];
                                countcolor_in = ninein_bitmap32[y_32][31-x_32];
                            end 
                            endcase
                        end
                        end
                    endcase
                end


                // 카운트다운용 카운터 
                if (clk_counter == 25_000_000 - 1) begin
                    clk_counter_next = 0;  // 카운터 초기화
                    if (countdown > 0) begin
                        countdown_next = countdown - 1;  // 카운트다운 감소
                    end else begin
                        countdown_next = 0;  // 카운트다운이 0이 되면 유지
                    end
                end else begin
                    clk_counter_next = clk_counter + 1;  // 카운터 증가
                end


                if (countdown == 0) begin
                    countdown_done_next = 1;  // 카운트다운 완료 신호
                    q_display_done_next = 0;
                    state_next = WIN_LOSE;        
                end 
            end







        /************************************LEVEL2-1******************************************/
        /************************************LEVEL2-1******************************************/
        /************************************LEVEL2-1******************************************/
        /************************************LEVEL2-1******************************************/
        /************************************LEVEL2-1******************************************/
        /************************************LEVEL2-1******************************************/
        /************************************LEVEL2-1******************************************/
        /************************************LEVEL2-1******************************************/
        /************************************LEVEL2-1******************************************/
        /************************************LEVEL2-1******************************************/
            LEVEL2_1: // 깜빡 + 한번에 2개 
            begin
                // blink counter
                game_done_next = 1;
                led_next = 4'b0011;
                if (clk_counter_blink == 2_500_000 - 1) begin
                    clk_counter_blink_next = 0;  // 카운터 초기화
                    if (blink_count == 49) begin
                        blink_count_next = 0;
                    end else begin
                        blink_count_next = blink_count + 1;
                    end
                end else begin
                    clk_counter_blink_next = clk_counter_blink + 1;  // 카운터 증가
                end



                // 게임 색깔 표시 (2개) (y= 80~200, x= 150 ~ 270) , (y= 80~200, x= 370 ~ 490)  
                if ((x_pixel < 270 && x_pixel >= 150) && (y_pixel < 200 && y_pixel >= 80)) begin         
                    if (blink_count == 1) begin
                        case (question[1:0])
                            2'd0: {red_port, green_port, blue_port} = {4'h0, 4'h0, 4'h0}; //black 0 들어오면 검정색
                            2'd1: {red_port, green_port, blue_port} = {4'hf, 4'h0, 4'h0}; //red
                            2'd2: {red_port, green_port, blue_port} = {4'hf, 4'hf, 4'h0}; //yellow
                            2'd3: {red_port, green_port, blue_port} = {4'h0, 4'h0, 4'hf}; //blue
                        endcase    
                    end else begin
                        {red_port, green_port, blue_port} = {cam_r, cam_g, cam_b}; // 깜빡이지 않을떈 아무것도 표시 X
                    end
                end else if ((x_pixel < 490 && x_pixel >= 370) && (y_pixel < 200 && y_pixel >= 80)) begin         
                    if (blink_count == 1) begin
                        q_display_done_next = 1;
                        case (question[3:2])
                            2'd0: {red_port, green_port, blue_port} = {4'h0, 4'h0, 4'h0}; //black 0 들어오면 검정색
                            2'd1: {red_port, green_port, blue_port} = {4'hf, 4'h0, 4'h0}; //red
                            2'd2: {red_port, green_port, blue_port} = {4'hf, 4'hf, 4'h0}; //yellow
                            2'd3: {red_port, green_port, blue_port} = {4'h0, 4'h0, 4'hf}; //blue
                        endcase    
                    end else begin
                        {red_port, green_port, blue_port} = {cam_r, cam_g, cam_b}; // 깜빡이지 않을떈 아무것도 표시 X
                    end
                end 



                // 정답 제출할 영역 표시 (검정색) , (y= 280~400, x= 150 ~ 270), (y= 280~400, x= 370 ~ 490)  
                else if (((x_pixel < 270 && x_pixel >= 150) && (y_pixel == 280 || y_pixel == 400)) ||
                        ((x_pixel == 270 || x_pixel == 150) && (y_pixel >= 280 && y_pixel < 400))) begin
                    red_port   = 4'h0;  // Red
                    green_port = 4'h0;  // Green
                    blue_port  = 4'h0;  // Blue  
                end else if (((x_pixel < 490 && x_pixel >= 370) && (y_pixel == 280 || y_pixel == 400)) ||
                        ((x_pixel == 490 || x_pixel == 370) && (y_pixel >= 280 && y_pixel < 400))) begin
                    red_port   = 4'h0;  // Red
                    green_port = 4'h0;  // Green
                    blue_port  = 4'h0;  // Blue  
                end



                // LEVEL 2 - 1 표시 (y= 28~60, x= 210 ~ 436) 
                else if (y_pixel >= 28 && y_pixel < 60) begin
                    y_32 = y_pixel - 28;
                    case (x_pixel) inside
                        [210:241]: begin        // L
                            x_32 = x_pixel - (210);
                            font_out = Lout_bitmap32[y_32][31-x_32];
                            font_in = Lin_bitmap32[y_32][31-x_32];
                        end
                        [243:274]: begin        // E
                            x_32 = x_pixel - (243);
                            font_out = Eout_bitmap32[y_32][31-x_32];
                            font_in = Ein_bitmap32[y_32][31-x_32];
                        end
                        [276:307]: begin        // V
                            x_32 = x_pixel - (276);
                            font_out = Vout_bitmap32[y_32][31-x_32];
                            font_in = Vin_bitmap32[y_32][31-x_32];
                        end
                        [309:340]: begin        // E
                            x_32 = x_pixel - (309);
                            font_out = Eout_bitmap32[y_32][31-x_32];
                            font_in = Ein_bitmap32[y_32][31-x_32];
                        end
                        [342:373]: begin        // L
                            x_32 = x_pixel - (342);
                            font_out = Lout_bitmap32[y_32][31-x_32];
                            font_in = Lin_bitmap32[y_32][31-x_32];
                        end
                        [405:436]: begin        // 2
                            x_32 = x_pixel - (405);
                            font_out = twoout_bitmap32[y_32][31-x_32];
                            font_in = twoin_bitmap32[y_32][31-x_32];
                        end
                        [440:471]: begin        // -
                            x_32 = x_pixel - (440);
                            font_out = dashout_bitmap32[y_32][31-x_32];
                            font_in = dashin_bitmap32[y_32][31-x_32];
                        end
                        [475:506]: begin        // 1
                            x_32 = x_pixel - (475);
                            font_out = oneout_bitmap32[y_32][31-x_32];
                            font_in = onein_bitmap32[y_32][31-x_32];
                        end
                        [550:581]: begin       // countdown (y= 28~60, x=500~532 )
                            if (q_display_done) begin
                            x_32 = x_pixel - (550);
                            case (countdown)
                            4'd0: begin
                                font_out = zeroout_bitmap32[y_32][31-x_32];
                                countcolor_in = zeroin_bitmap32[y_32][31-x_32];
                            end 
                            4'd1: begin
                                font_out = oneout_bitmap32[y_32][31-x_32];
                                countcolor_in = onein_bitmap32[y_32][31-x_32];
                            end 
                            4'd2: begin
                                font_out = twoout_bitmap32[y_32][31-x_32];
                                countcolor_in = twoin_bitmap32[y_32][31-x_32];
                            end 
                            4'd3: begin
                                font_out = threeout_bitmap32[y_32][31-x_32];
                                countcolor_in = threein_bitmap32[y_32][31-x_32];
                            end 
                            4'd4: begin
                                font_out = fourout_bitmap32[y_32][31-x_32];
                                countcolor_in = fourin_bitmap32[y_32][31-x_32];
                            end 
                            4'd5: begin
                                font_out = fiveout_bitmap32[y_32][31-x_32];
                                countcolor_in = fivein_bitmap32[y_32][31-x_32];
                            end 
                            4'd6: begin
                                font_out = sixout_bitmap32[y_32][31-x_32];
                                countcolor_in = sixin_bitmap32[y_32][31-x_32];
                            end 
                            4'd7: begin
                                font_out = sevenout_bitmap32[y_32][31-x_32];
                                countcolor_in = sevenin_bitmap32[y_32][31-x_32];
                            end 
                            4'd8: begin
                                font_out = eightout_bitmap32[y_32][31-x_32];
                                countcolor_in = eightin_bitmap32[y_32][31-x_32];
                            end 
                            4'd9: begin
                                font_out = nineout_bitmap32[y_32][31-x_32];
                                countcolor_in = ninein_bitmap32[y_32][31-x_32];
                            end 
                            endcase
                            end
                        end
                    endcase
                end
                

                // 카운트 다운용 카운터 
                if (clk_counter == 25_000_000 - 1) begin
                    clk_counter_next = 0;  // 카운터 초기화
                    if (countdown > 0) begin
                        countdown_next = countdown - 1;  // 카운트다운 감소
                    end else begin
                        countdown_next = 0;  // 카운트다운이 0이 되면 유지
                    end
                end else begin
                    clk_counter_next = clk_counter + 1;  // 카운터 증가
                end

                if (countdown == 0) begin
                    countdown_done_next = 1;  // 카운트다운 완료 신호
                    q_display_done_next = 0;
                    state_next = WIN_LOSE;
                end 
            end

        LEVEL2_2: // 깜빡 + 한번에 3개 
            begin
                // blink counter
                game_done_next = 1;
                led_next = 4'b0011;
                if (clk_counter_blink == 2_500_000 - 1) begin
                    clk_counter_blink_next = 0;  // 카운터 초기화
                    if (blink_count == 49) begin
                        blink_count_next = 0;
                    end else begin
                        blink_count_next = blink_count + 1;
                    end
                end else begin
                    clk_counter_blink_next = clk_counter_blink + 1;  // 카운터 증가
                end



                // 게임 색깔 표시 (3개) (y= 80~200, x= 70 ~ 190) , (y= 80~200, x= 260 ~ 380) , (y= 80~200, x= 450 ~ 570) 
                if ((x_pixel < 190 && x_pixel >= 70) && (y_pixel < 200 && y_pixel >= 80)) begin         
                    if (blink_count == 1) begin
                        q_display_done_next = 1;
                        case (question[1:0])
                            2'd0: {red_port, green_port, blue_port} = {4'h0, 4'h0, 4'h0}; //black 0 들어오면 검정색
                            2'd1: {red_port, green_port, blue_port} = {4'hf, 4'h0, 4'h0}; //red
                            2'd2: {red_port, green_port, blue_port} = {4'hf, 4'hf, 4'h0}; //yellow
                            2'd3: {red_port, green_port, blue_port} = {4'h0, 4'h0, 4'hf}; //blue
                        endcase    
                    end else begin
                        {red_port, green_port, blue_port} = {cam_r, cam_g, cam_b}; // 깜빡이지 않을떈 아무것도 표시 X
                    end
                end else if ((x_pixel < 380 && x_pixel >= 260) && (y_pixel < 200 && y_pixel >= 80)) begin         
                    if (blink_count == 1) begin
                        case (question[3:2])
                            2'd0: {red_port, green_port, blue_port} = {4'h0, 4'h0, 4'h0}; //black 0 들어오면 검정색
                            2'd1: {red_port, green_port, blue_port} = {4'hf, 4'h0, 4'h0}; //red
                            2'd2: {red_port, green_port, blue_port} = {4'hf, 4'hf, 4'h0}; //yellow
                            2'd3: {red_port, green_port, blue_port} = {4'h0, 4'h0, 4'hf}; //blue
                        endcase    
                    end else begin
                        {red_port, green_port, blue_port} = {cam_r, cam_g, cam_b}; // 깜빡이지 않을떈 아무것도 표시 X
                    end
                end else if ((x_pixel < 570 && x_pixel >= 450) && (y_pixel < 200 && y_pixel >= 80)) begin         
                    if (blink_count == 1) begin
                        case (question[5:4])
                            2'd0: {red_port, green_port, blue_port} = {4'h0, 4'h0, 4'h0}; //black 0 들어오면 검정색
                            2'd1: {red_port, green_port, blue_port} = {4'hf, 4'h0, 4'h0}; //red
                            2'd2: {red_port, green_port, blue_port} = {4'hf, 4'hf, 4'h0}; //yellow
                            2'd3: {red_port, green_port, blue_port} = {4'h0, 4'h0, 4'hf}; //blue
                        endcase    
                    end else begin
                        {red_port, green_port, blue_port} = {cam_r, cam_g, cam_b}; // 깜빡이지 않을떈 아무것도 표시 X
                    end
                end 



                // 정답 제출할 영역 표시 (y= 280~400, x= 70 ~ 190), (y= 280~400, x= 260 ~ 380) , (y= 280~400, x= 450 ~ 570)  
                else if (((x_pixel < 190 && x_pixel >= 70) && (y_pixel == 280 || y_pixel == 400)) ||
                        ((x_pixel == 190 || x_pixel == 70) && (y_pixel >= 280 && y_pixel < 400))) begin
                    red_port   = 4'h0;  
                    green_port = 4'h0;  
                    blue_port  = 4'h0;  // -> black 
                end else if (((x_pixel < 380 && x_pixel >= 260) && (y_pixel == 280 || y_pixel == 400)) ||
                        ((x_pixel == 380 || x_pixel == 260) && (y_pixel >= 280 && y_pixel < 400))) begin
                    red_port   = 4'h0;  
                    green_port = 4'h0;  
                    blue_port  = 4'h0;  // -> black  
                end else if (((x_pixel < 570 && x_pixel >= 450) && (y_pixel == 280 || y_pixel == 400)) ||
                        ((x_pixel == 570 || x_pixel == 450) && (y_pixel >= 280 && y_pixel < 400))) begin
                    red_port   = 4'h0;  
                    green_port = 4'h0;  
                    blue_port  = 4'h0;  // -> black  
                end 



                // LEVEL 2-2 표시 (y= 28~60, x= 210 ~ 436) 
                else if (y_pixel >= 28 && y_pixel < 60) begin
                    y_32 = y_pixel - 28;
                    case (x_pixel) inside
                        [210:241]: begin        // L
                            x_32 = x_pixel - (210);
                            font_out = Lout_bitmap32[y_32][31-x_32];
                            font_in = Lin_bitmap32[y_32][31-x_32];
                        end
                        [243:274]: begin        // E
                            x_32 = x_pixel - (243);
                            font_out = Eout_bitmap32[y_32][31-x_32];
                            font_in = Ein_bitmap32[y_32][31-x_32];
                        end
                        [276:307]: begin        // V
                            x_32 = x_pixel - (276);
                            font_out = Vout_bitmap32[y_32][31-x_32];
                            font_in = Vin_bitmap32[y_32][31-x_32];
                        end
                        [309:340]: begin        // E
                            x_32 = x_pixel - (309);
                            font_out = Eout_bitmap32[y_32][31-x_32];
                            font_in = Ein_bitmap32[y_32][31-x_32];
                        end
                        [342:373]: begin        // L
                            x_32 = x_pixel - (342);
                            font_out = Lout_bitmap32[y_32][31-x_32];
                            font_in = Lin_bitmap32[y_32][31-x_32];
                        end
                        [405:436]: begin        // 2
                            x_32 = x_pixel - (405);
                            font_out = twoout_bitmap32[y_32][31-x_32];
                            font_in = twoin_bitmap32[y_32][31-x_32];
                        end
                        [440:471]: begin        // -
                            x_32 = x_pixel - (440);
                            font_out = dashout_bitmap32[y_32][31-x_32];
                            font_in = dashin_bitmap32[y_32][31-x_32];
                        end
                        [475:506]: begin        // 2
                            x_32 = x_pixel - (475);
                            font_out = twoout_bitmap32[y_32][31-x_32];
                            font_in = twoin_bitmap32[y_32][31-x_32];
                        end
                        [550:581]: begin       // countdown (y= 28~60, x=500~532 )
                            if (q_display_done) begin
                            x_32 = x_pixel - (550);
                            case (countdown)
                            4'd0: begin
                                font_out = zeroout_bitmap32[y_32][31-x_32];
                                countcolor_in = zeroin_bitmap32[y_32][31-x_32];
                            end 
                            4'd1: begin
                                font_out = oneout_bitmap32[y_32][31-x_32];
                                countcolor_in = onein_bitmap32[y_32][31-x_32];
                            end 
                            4'd2: begin
                                font_out = twoout_bitmap32[y_32][31-x_32];
                                countcolor_in = twoin_bitmap32[y_32][31-x_32];
                            end 
                            4'd3: begin
                                font_out = threeout_bitmap32[y_32][31-x_32];
                                countcolor_in = threein_bitmap32[y_32][31-x_32];
                            end 
                            4'd4: begin
                                font_out = fourout_bitmap32[y_32][31-x_32];
                                countcolor_in = fourin_bitmap32[y_32][31-x_32];
                            end 
                            4'd5: begin
                                font_out = fiveout_bitmap32[y_32][31-x_32];
                                countcolor_in = fivein_bitmap32[y_32][31-x_32];
                            end 
                            4'd6: begin
                                font_out = sixout_bitmap32[y_32][31-x_32];
                                countcolor_in = sixin_bitmap32[y_32][31-x_32];
                            end 
                            4'd7: begin
                                font_out = sevenout_bitmap32[y_32][31-x_32];
                                countcolor_in = sevenin_bitmap32[y_32][31-x_32];
                            end 
                            4'd8: begin
                                font_out = eightout_bitmap32[y_32][31-x_32];
                                countcolor_in = eightin_bitmap32[y_32][31-x_32];
                            end 
                            4'd9: begin
                                font_out = nineout_bitmap32[y_32][31-x_32];
                                countcolor_in = ninein_bitmap32[y_32][31-x_32];
                            end 
                            endcase
                            end
                        end
                    endcase
                end
                

                // 카운트 다운용 카운터 
                if (clk_counter == 25_000_000 - 1) begin
                    clk_counter_next = 0;  // 카운터 초기화
                    if (countdown > 0) begin
                        countdown_next = countdown - 1;  // 카운트다운 감소
                    end else begin
                        countdown_next = 0;  // 카운트다운이 0이 되면 유지
                    end
                end else begin
                    clk_counter_next = clk_counter + 1;  // 카운터 증가
                end

                if (countdown == 0) begin
                    countdown_done_next = 1;  // 카운트다운 완료 신호
                    q_display_done_next = 0;
                    state_next = WIN_LOSE;
                end 
            end

            LEVEL2_3: // 깜빡 + 한번에 4개 
            begin
                // blink counter
                game_done_next = 1;
                led_next = 4'b0011;
                if (clk_counter_blink == 2_500_000 - 1) begin
                    clk_counter_blink_next = 0;  // 카운터 초기화
                    if (blink_count == 49) begin
                        blink_count_next = 0;
                    end else begin
                        blink_count_next = blink_count + 1;
                    end
                end else begin
                    clk_counter_blink_next = clk_counter_blink + 1;  // 카운터 증가
                end



                // 게임 색깔 표시 (4개) (y= 80~200, x= 32 ~ 152) , (y= 80~200, x= 184 ~ 304) , (y= 80~200, x= 336 ~ 456) , (y= 80~200, x= 488 ~ 608) 
                if ((x_pixel < 152 && x_pixel >= 32) && (y_pixel < 200 && y_pixel >= 80)) begin         
                    if (blink_count == 1) begin
                        q_display_done_next = 1;
                        case (question[1:0])
                            2'd0: {red_port, green_port, blue_port} = {4'h0, 4'h0, 4'h0}; //black 0 들어오면 검정색
                            2'd1: {red_port, green_port, blue_port} = {4'hf, 4'h0, 4'h0}; //red
                            2'd2: {red_port, green_port, blue_port} = {4'hf, 4'hf, 4'h0}; //yellow
                            2'd3: {red_port, green_port, blue_port} = {4'h0, 4'h0, 4'hf}; //blue
                        endcase    
                    end else begin
                        {red_port, green_port, blue_port} = {cam_r, cam_g, cam_b}; // 깜빡이지 않을떈 아무것도 표시 X
                    end
                end else if ((x_pixel < 304 && x_pixel >= 184) && (y_pixel < 200 && y_pixel >= 80)) begin         
                    if (blink_count == 1) begin
                        case (question[3:2])
                            2'd0: {red_port, green_port, blue_port} = {4'h0, 4'h0, 4'h0}; //black 0 들어오면 검정색
                            2'd1: {red_port, green_port, blue_port} = {4'hf, 4'h0, 4'h0}; //red
                            2'd2: {red_port, green_port, blue_port} = {4'hf, 4'hf, 4'h0}; //yellow
                            2'd3: {red_port, green_port, blue_port} = {4'h0, 4'h0, 4'hf}; //blue
                        endcase    
                    end else begin
                        {red_port, green_port, blue_port} = {cam_r, cam_g, cam_b}; // 깜빡이지 않을떈 아무것도 표시 X
                    end
                end else if ((x_pixel < 456 && x_pixel >= 336) && (y_pixel < 200 && y_pixel >= 80)) begin         
                    if (blink_count == 1) begin
                        case (question[5:4])
                            2'd0: {red_port, green_port, blue_port} = {4'h0, 4'h0, 4'h0}; //black 0 들어오면 검정색
                            2'd1: {red_port, green_port, blue_port} = {4'hf, 4'h0, 4'h0}; //red
                            2'd2: {red_port, green_port, blue_port} = {4'hf, 4'hf, 4'h0}; //yellow
                            2'd3: {red_port, green_port, blue_port} = {4'h0, 4'h0, 4'hf}; //blue
                        endcase    
                    end else begin
                        {red_port, green_port, blue_port} = {cam_r, cam_g, cam_b}; // 깜빡이지 않을떈 아무것도 표시 X
                    end
                end else if ((x_pixel < 608 && x_pixel >= 488) && (y_pixel < 200 && y_pixel >= 80)) begin         
                    if (blink_count == 1) begin
                        case (question[7:6])
                            2'd0: {red_port, green_port, blue_port} = {4'h0, 4'h0, 4'h0}; //black 0 들어오면 검정색
                            2'd1: {red_port, green_port, blue_port} = {4'hf, 4'h0, 4'h0}; //red
                            2'd2: {red_port, green_port, blue_port} = {4'hf, 4'hf, 4'h0}; //yellow
                            2'd3: {red_port, green_port, blue_port} = {4'h0, 4'h0, 4'hf}; //blue
                        endcase    
                    end else begin
                        {red_port, green_port, blue_port} = {cam_r, cam_g, cam_b}; // 깜빡이지 않을떈 아무것도 표시 X
                    end
                end 



                // 정답 제출할 영역 표시 (y= 280~400, x= 32 ~ 152), (y= 280~400, x= 184 ~ 304) , (y= 280~400, x= 336 ~ 456)  , (y= 280~400, x= 488 ~ 608)  
                else if (((x_pixel < 152 && x_pixel >= 32) && (y_pixel == 280 || y_pixel == 400)) ||
                        ((x_pixel == 152 || x_pixel == 32) && (y_pixel >= 280 && y_pixel < 400))) begin
                    red_port   = 4'h0;  
                    green_port = 4'h0;  
                    blue_port  = 4'h0;  // -> black 
                end else if (((x_pixel < 304 && x_pixel >= 184) && (y_pixel == 280 || y_pixel == 400)) ||
                            ((x_pixel == 304 || x_pixel == 184) && (y_pixel >= 280 && y_pixel < 400))) begin
                    red_port   = 4'h0;  
                    green_port = 4'h0;  
                    blue_port  = 4'h0;  // -> black  
                end else if (((x_pixel < 456 && x_pixel >= 336) && (y_pixel == 280 || y_pixel == 400)) ||
                            ((x_pixel == 456 || x_pixel == 336) && (y_pixel >= 280 && y_pixel < 400))) begin
                    red_port   = 4'h0;  
                    green_port = 4'h0;  
                    blue_port  = 4'h0;  // -> black  
                end else if (((x_pixel < 608 && x_pixel >= 488) && (y_pixel == 280 || y_pixel == 400)) ||
                            ((x_pixel == 608 || x_pixel == 488) && (y_pixel >= 280 && y_pixel < 400))) begin
                    red_port   = 4'h0;  
                    green_port = 4'h0;  
                    blue_port  = 4'h0;  // -> black  
                end 



                // LEVEL 2-3 표시 (y= 28~60, x= 210 ~ 436) 
                else if (y_pixel >= 28 && y_pixel < 60) begin
                    y_32 = y_pixel - 28;
                    case (x_pixel) inside
                        [210:241]: begin        // L
                            x_32 = x_pixel - (210);
                            font_out = Lout_bitmap32[y_32][31-x_32];
                            font_in = Lin_bitmap32[y_32][31-x_32];
                        end
                        [243:274]: begin        // E
                            x_32 = x_pixel - (243);
                            font_out = Eout_bitmap32[y_32][31-x_32];
                            font_in = Ein_bitmap32[y_32][31-x_32];
                        end
                        [276:307]: begin        // V
                            x_32 = x_pixel - (276);
                            font_out = Vout_bitmap32[y_32][31-x_32];
                            font_in = Vin_bitmap32[y_32][31-x_32];
                        end
                        [309:340]: begin        // E
                            x_32 = x_pixel - (309);
                            font_out = Eout_bitmap32[y_32][31-x_32];
                            font_in = Ein_bitmap32[y_32][31-x_32];
                        end
                        [342:373]: begin        // L
                            x_32 = x_pixel - (342);
                            font_out = Lout_bitmap32[y_32][31-x_32];
                            font_in = Lin_bitmap32[y_32][31-x_32];
                        end
                        [405:436]: begin        // 2
                            x_32 = x_pixel - (405);
                            font_out = twoout_bitmap32[y_32][31-x_32];
                            font_in = twoin_bitmap32[y_32][31-x_32];
                        end
                        [440:471]: begin        // -
                            x_32 = x_pixel - (440);
                            font_out = dashout_bitmap32[y_32][31-x_32];
                            font_in = dashin_bitmap32[y_32][31-x_32];
                        end
                        [475:506]: begin        // 3
                            x_32 = x_pixel - (475);
                            font_out = threeout_bitmap32[y_32][31-x_32];
                            font_in = threein_bitmap32[y_32][31-x_32];
                        end
                        [550:581]: begin       // countdown (y= 28~60, x=500~532 )
                            if (q_display_done) begin
                            x_32 = x_pixel - (550);
                            case (countdown)
                            4'd0: begin
                                font_out = zeroout_bitmap32[y_32][31-x_32];
                                countcolor_in = zeroin_bitmap32[y_32][31-x_32];
                            end 
                            4'd1: begin
                                font_out = oneout_bitmap32[y_32][31-x_32];
                                countcolor_in = onein_bitmap32[y_32][31-x_32];
                            end 
                            4'd2: begin
                                font_out = twoout_bitmap32[y_32][31-x_32];
                                countcolor_in = twoin_bitmap32[y_32][31-x_32];
                            end 
                            4'd3: begin
                                font_out = threeout_bitmap32[y_32][31-x_32];
                                countcolor_in = threein_bitmap32[y_32][31-x_32];
                            end 
                            4'd4: begin
                                font_out = fourout_bitmap32[y_32][31-x_32];
                                countcolor_in = fourin_bitmap32[y_32][31-x_32];
                            end 
                            4'd5: begin
                                font_out = fiveout_bitmap32[y_32][31-x_32];
                                countcolor_in = fivein_bitmap32[y_32][31-x_32];
                            end 
                            4'd6: begin
                                font_out = sixout_bitmap32[y_32][31-x_32];
                                countcolor_in = sixin_bitmap32[y_32][31-x_32];
                            end 
                            4'd7: begin
                                font_out = sevenout_bitmap32[y_32][31-x_32];
                                countcolor_in = sevenin_bitmap32[y_32][31-x_32];
                            end 
                            4'd8: begin
                                font_out = eightout_bitmap32[y_32][31-x_32];
                                countcolor_in = eightin_bitmap32[y_32][31-x_32];
                            end 
                            4'd9: begin
                                font_out = nineout_bitmap32[y_32][31-x_32];
                                countcolor_in = ninein_bitmap32[y_32][31-x_32];
                            end 
                            endcase
                            end
                        end
                    endcase
                end
                

                // 카운트 다운용 카운터 
                if (clk_counter == 25_000_000 - 1) begin
                    clk_counter_next = 0;  // 카운터 초기화
                    if (countdown > 0) begin
                        countdown_next = countdown - 1;  // 카운트다운 감소
                    end else begin
                        countdown_next = 0;  // 카운트다운이 0이 되면 유지
                    end
                end else begin
                    clk_counter_next = clk_counter + 1;  // 카운터 증가
                end

                if (countdown == 0) begin
                    countdown_done_next = 1;  // 카운트다운 완료 신호
                    q_display_done_next = 0;
                    state_next = WIN_LOSE;
                end 
            end


        /************************************LEVEL3******************************************/
        /************************************LEVEL3******************************************/
        /************************************LEVEL3******************************************/
        /************************************LEVEL3******************************************/
        /************************************LEVEL3******************************************/
        /************************************LEVEL3******************************************/
        /************************************LEVEL3******************************************/
        /************************************LEVEL3******************************************/
        /************************************LEVEL3******************************************/
        /************************************LEVEL3******************************************/
            LEVEL3_1: // Blink + 글자 4개 (글자와 색깔 다르게)
            begin
                // blink counter
                led_next = 4'b0100;
                if (clk_counter_blink == 2_500_000 - 1) begin
                    clk_counter_blink_next = 0;  // 카운터 초기화
                    if (blink_count == 49) begin
                        blink_count_next = 0;
                    end else begin
                        blink_count_next = blink_count + 1;
                    end
                end else begin
                    clk_counter_blink_next = clk_counter_blink + 1;  // 카운터 증가
                end



                 // 게임 색깔 표시 (4개) (y= 80~200, x= 32 ~ 152) , (y= 80~200, x= 184 ~ 304) , (y= 80~200, x= 336 ~ 456) , (y= 80~200, x= 488 ~ 608) 
                if (y_pixel >= 124 && y_pixel < 156) begin
                        y_32 = y_pixel - 124;
                        q_display_done_next = 1;
                        case (x_pixel) inside
                        [150:270]:begin
                            case (question[1:0])
                                2'd0: {red_port, green_port, blue_port} = {4'h0, 4'h0, 4'h0}; //black 0 들어오면 검정색
                                2'd1: begin     //RED
                                        case (x_pixel) inside
                                            [154:185]: begin        // R
                                                x_32 = x_pixel - (154);
                                                font_out = Rout_bitmap32[y_32][31-x_32];
                                                Y_in = Rin_bitmap32[y_32][31-x_32];
                                            end
                                            [194:225]: begin        // E
                                                x_32 = x_pixel - (194);
                                                font_out = Eout_bitmap32[y_32][31-x_32];
                                                Y_in = Ein_bitmap32[y_32][31-x_32];
                                            end
                                            [234:265]: begin        // D
                                                x_32 = x_pixel - (234);
                                                font_out = Dout_bitmap32[y_32][31-x_32];
                                                Y_in = Din_bitmap32[y_32][31-x_32];
                                            end
                                        endcase
                                end
                                2'd2: case (x_pixel) inside
                                            [154:185]: begin        // Y
                                                x_32 = x_pixel - (154);
                                                font_out = Yout_bitmap32[y_32][31-x_32];
                                                B_in = Yin_bitmap32[y_32][31-x_32];
                                            end
                                            [194:225]: begin        // E
                                                x_32 = x_pixel - (194);
                                                font_out = Eout_bitmap32[y_32][31-x_32];
                                                B_in = Ein_bitmap32[y_32][31-x_32];
                                            end
                                            [234:265]: begin      // L
                                                x_32 = x_pixel - (234);
                                                font_out = Lout_bitmap32[y_32][31-x_32];
                                                B_in = Lin_bitmap32[y_32][31-x_32];
                                            end
                                        endcase //yellow
                                2'd3: case (x_pixel) inside
                                            [154:185]: begin        // B
                                                x_32 = x_pixel - (154);
                                                font_out = Bout_bitmap32[y_32][31-x_32];
                                                G_in = Bin_bitmap32[y_32][31-x_32];
                                            end
                                            [194:225]: begin        // L
                                                x_32 = x_pixel - (194);
                                                font_out = Lout_bitmap32[y_32][31-x_32];
                                                G_in = Lin_bitmap32[y_32][31-x_32];
                                            end
                                            [234:265]: begin      // U
                                                x_32 = x_pixel - (234);
                                                font_out = Uout_bitmap32[y_32][31-x_32];
                                                G_in = Uin_bitmap32[y_32][31-x_32];
                                            end
                                        endcase //blue
                            endcase
                        end
                        [370:490]: begin
                            case (question[3:2])
                                2'd0: {red_port, green_port, blue_port} = {4'h0, 4'h0, 4'h0}; //black 0 들어오면 검정색
                                2'd1: begin     //YELLOW
                                        case (x_pixel) inside
                                            [374:405]: begin        // R
                                                x_32 = x_pixel - (374);
                                                font_out = Rout_bitmap32[y_32][31-x_32];
                                                B_in = Rin_bitmap32[y_32][31-x_32];
                                            end
                                            [414:445]: begin        // E
                                                x_32 = x_pixel - (414);
                                                font_out = Eout_bitmap32[y_32][31-x_32];
                                                B_in = Ein_bitmap32[y_32][31-x_32];
                                            end
                                            [454:485]: begin        // D
                                                x_32 = x_pixel - (454);
                                                font_out = Dout_bitmap32[y_32][31-x_32];
                                                B_in = Din_bitmap32[y_32][31-x_32];
                                            end
                                        endcase
                                end //red
                                2'd2: begin     //YELLOW
                                        case (x_pixel) inside
                                            [374:405]: begin        // Y
                                                x_32 = x_pixel - (374);
                                                font_out = Yout_bitmap32[y_32][31-x_32];
                                                R_in = Yin_bitmap32[y_32][31-x_32];
                                            end
                                            [414:445]: begin        // E
                                                x_32 = x_pixel - (414);
                                                font_out = Eout_bitmap32[y_32][31-x_32];
                                                R_in = Ein_bitmap32[y_32][31-x_32];
                                            end
                                            [454:485]: begin        // L
                                                x_32 = x_pixel - (454);
                                                font_out = Lout_bitmap32[y_32][31-x_32];
                                                R_in = Lin_bitmap32[y_32][31-x_32];
                                            end
                                        endcase
                                end
                                2'd3: begin     //YELLOW
                                        case (x_pixel) inside
                                            [374:405]: begin        // B
                                                x_32 = x_pixel - (374);
                                                font_out = Bout_bitmap32[y_32][31-x_32];
                                                P_in = Bin_bitmap32[y_32][31-x_32];
                                            end
                                            [414:445]: begin        // L
                                                x_32 = x_pixel - (414);
                                                font_out = Lout_bitmap32[y_32][31-x_32];
                                                P_in = Lin_bitmap32[y_32][31-x_32];
                                            end
                                            [454:485]: begin        // U
                                                x_32 = x_pixel - (454);
                                                font_out = Uout_bitmap32[y_32][31-x_32];
                                                P_in = Uin_bitmap32[y_32][31-x_32];
                                            end
                                        endcase
                                end //blue
                            endcase
                        end
                        default: {red_port, green_port, blue_port} = {cam_r, cam_g, cam_b};
                        endcase 
                    end 
                 
                


                // 정답 제출할 영역 표시 (y= 280~400, x= 32 ~ 152), (y= 280~400, x= 184 ~ 304) , (y= 280~400, x= 336 ~ 456)  , (y= 280~400, x= 488 ~ 608)  
                else if (((x_pixel < 270 && x_pixel >= 150) && (y_pixel == 280 || y_pixel == 400)) ||
                        ((x_pixel == 270 || x_pixel == 150) && (y_pixel >= 280 && y_pixel < 400))) begin
                    red_port   = 4'h0;  
                    green_port = 4'h0;  
                    blue_port  = 4'h0;  // -> black 
                end else if (((x_pixel < 490 && x_pixel >= 370) && (y_pixel == 280 || y_pixel == 400)) ||
                            ((x_pixel == 490 || x_pixel == 370) && (y_pixel >= 280 && y_pixel < 400))) begin
                    red_port   = 4'h0;  
                    green_port = 4'h0;  
                    blue_port  = 4'h0;  // -> black  
                end


                // LEVEL 3 표시 (y= 28~60, x= 210 ~ 436) 
                else if (y_pixel >= 28 && y_pixel < 60) begin
                    y_32 = y_pixel - 28;
                    case (x_pixel) inside
                        [210:241]: begin        // L
                            x_32 = x_pixel - (210);
                            font_out = Lout_bitmap32[y_32][31-x_32];
                            font_in = Lin_bitmap32[y_32][31-x_32];
                        end
                        [243:274]: begin        // E
                            x_32 = x_pixel - (243);
                            font_out = Eout_bitmap32[y_32][31-x_32];
                            font_in = Ein_bitmap32[y_32][31-x_32];
                        end
                        [276:307]: begin        // V
                            x_32 = x_pixel - (276);
                            font_out = Vout_bitmap32[y_32][31-x_32];
                            font_in = Vin_bitmap32[y_32][31-x_32];
                        end
                        [309:340]: begin        // E
                            x_32 = x_pixel - (309);
                            font_out = Eout_bitmap32[y_32][31-x_32];
                            font_in = Ein_bitmap32[y_32][31-x_32];
                        end
                        [342:373]: begin        // L
                            x_32 = x_pixel - (342);
                            font_out = Lout_bitmap32[y_32][31-x_32];
                            font_in = Lin_bitmap32[y_32][31-x_32];
                        end
                        [405:436]: begin        // 3
                            x_32 = x_pixel - (405);
                            font_out = threeout_bitmap32[y_32][31-x_32];
                            font_in = threein_bitmap32[y_32][31-x_32];
                        end
                        [440:471]: begin        // -
                            x_32 = x_pixel - (440);
                            font_out = dashout_bitmap32[y_32][31-x_32];
                            font_in = dashin_bitmap32[y_32][31-x_32];
                        end
                        [475:506]: begin        // 1
                            x_32 = x_pixel - (475);
                            font_out = oneout_bitmap32[y_32][31-x_32];
                            font_in = onein_bitmap32[y_32][31-x_32];
                        end
                        [550:581]: begin       // countdown (y= 28~60, x=500~532 )
                        if (q_display_done) begin
                            x_32 = x_pixel - (550);
                            case (countdown)
                            4'd0: begin
                                font_out = zeroout_bitmap32[y_32][31-x_32];
                                countcolor_in = zeroin_bitmap32[y_32][31-x_32];
                            end 
                            4'd1: begin
                                font_out = oneout_bitmap32[y_32][31-x_32];
                                countcolor_in = onein_bitmap32[y_32][31-x_32];
                            end 
                            4'd2: begin
                                font_out = twoout_bitmap32[y_32][31-x_32];
                                countcolor_in = twoin_bitmap32[y_32][31-x_32];
                            end 
                            4'd3: begin
                                font_out = threeout_bitmap32[y_32][31-x_32];
                                countcolor_in = threein_bitmap32[y_32][31-x_32];
                            end 
                            4'd4: begin
                                font_out = fourout_bitmap32[y_32][31-x_32];
                                countcolor_in = fourin_bitmap32[y_32][31-x_32];
                            end 
                            4'd5: begin
                                font_out = fiveout_bitmap32[y_32][31-x_32];
                                countcolor_in = fivein_bitmap32[y_32][31-x_32];
                            end 
                            4'd6: begin
                                font_out = sixout_bitmap32[y_32][31-x_32];
                                countcolor_in = sixin_bitmap32[y_32][31-x_32];
                            end 
                            4'd7: begin
                                font_out = sevenout_bitmap32[y_32][31-x_32];
                                countcolor_in = sevenin_bitmap32[y_32][31-x_32];
                            end 
                            4'd8: begin
                                font_out = eightout_bitmap32[y_32][31-x_32];
                                countcolor_in = eightin_bitmap32[y_32][31-x_32];
                            end 
                            4'd9: begin
                                font_out = nineout_bitmap32[y_32][31-x_32];
                                countcolor_in = ninein_bitmap32[y_32][31-x_32];
                            end 
                            endcase
                        end
                        end
                    endcase
                end
                

                // 카운트 다운용 카운터 
                if (clk_counter == 25_000_000 - 1) begin
                    clk_counter_next = 0;  // 카운터 초기화
                    if (countdown > 0) begin
                        countdown_next = countdown - 1;  // 카운트다운 감소
                    end else begin
                        countdown_next = 0;  // 카운트다운이 0이 되면 유지
                    end
                end else begin
                    clk_counter_next = clk_counter + 1;  // 카운터 증가
                end

                if (countdown == 0) begin
                    countdown_done_next = 1;  // 카운트다운 완료 신호
                    q_display_done_next = 0;
                    // win 
                    state_next = WIN_LOSE;
                end 
            end
            
            LEVEL3_2: // Blink + 글자 4개 (글자와 색깔 다르게)
            begin
                // blink counter
                led_next = 4'b0100;
                if (clk_counter_blink == 2_500_000 - 1) begin
                    clk_counter_blink_next = 0;  // 카운터 초기화
                    if (blink_count == 49) begin
                        blink_count_next = 0;
                    end else begin
                        blink_count_next = blink_count + 1;
                    end
                end else begin
                    clk_counter_blink_next = clk_counter_blink + 1;  // 카운터 증가
                end



                 // 게임 색깔 표시 (4개) (y= 80~200, x= 32 ~ 152) , (y= 80~200, x= 184 ~ 304) , (y= 80~200, x= 336 ~ 456) , (y= 80~200, x= 488 ~ 608) 
                if (y_pixel >= 124 && y_pixel < 156) begin
                        y_32 = y_pixel - 124;
                        q_display_done_next = 1;
                        case (x_pixel) inside
                        [70:190]:begin
                            case (question[1:0])
                                2'd0: {red_port, green_port, blue_port} = {4'h0, 4'h0, 4'h0}; //black 0 들어오면 검정색
                                2'd1: begin     //RED
                                        case (x_pixel) inside
                                            [74:105]: begin        // R
                                                x_32 = x_pixel - (74);
                                                font_out = Rout_bitmap32[y_32][31-x_32];
                                                G_in = Rin_bitmap32[y_32][31-x_32];
                                            end
                                            [114:145]: begin        // E
                                                x_32 = x_pixel - (114);
                                                font_out = Eout_bitmap32[y_32][31-x_32];
                                                G_in = Ein_bitmap32[y_32][31-x_32];
                                            end
                                            [154:185]: begin        // D
                                                x_32 = x_pixel - (154);
                                                font_out = Dout_bitmap32[y_32][31-x_32];
                                                G_in = Din_bitmap32[y_32][31-x_32];
                                            end
                                        endcase
                                end
                                2'd2: case (x_pixel) inside
                                            [74:105]: begin        // Y
                                                x_32 = x_pixel - (74);
                                                font_out = Yout_bitmap32[y_32][31-x_32];
                                                P_in = Yin_bitmap32[y_32][31-x_32];
                                            end
                                            [114:145]: begin        // E
                                                x_32 = x_pixel - (114);
                                                font_out = Eout_bitmap32[y_32][31-x_32];
                                                P_in = Ein_bitmap32[y_32][31-x_32];
                                            end
                                            [154:185]: begin      // L
                                                x_32 = x_pixel - (154);
                                                font_out = Lout_bitmap32[y_32][31-x_32];
                                                P_in = Lin_bitmap32[y_32][31-x_32];
                                            end
                                        endcase //yellow
                                2'd3: case (x_pixel) inside
                                            [74:105]: begin        // B
                                                x_32 = x_pixel - (74);
                                                font_out = Bout_bitmap32[y_32][31-x_32];
                                                Y_in = Bin_bitmap32[y_32][31-x_32];
                                            end
                                            [114:145]: begin        // L
                                                x_32 = x_pixel - (114);
                                                font_out = Lout_bitmap32[y_32][31-x_32];
                                                Y_in = Lin_bitmap32[y_32][31-x_32];
                                            end
                                            [154:185]: begin      // U
                                                x_32 = x_pixel - (154);
                                                font_out = Uout_bitmap32[y_32][31-x_32];
                                                Y_in = Uin_bitmap32[y_32][31-x_32];
                                            end
                                        endcase //blue
                            endcase
                        end
                        [260:380]: begin
                            case (question[3:2])
                                2'd0: {red_port, green_port, blue_port} = {4'h0, 4'h0, 4'h0}; //black 0 들어오면 검정색
                                2'd1: begin     //YELLOW
                                        case (x_pixel) inside
                                            [264:295]: begin        // R
                                                x_32 = x_pixel - (264);
                                                font_out = Rout_bitmap32[y_32][31-x_32];
                                                Y_in = Rin_bitmap32[y_32][31-x_32];
                                            end
                                            [304:335]: begin        // E
                                                x_32 = x_pixel - (304);
                                                font_out = Eout_bitmap32[y_32][31-x_32];
                                                Y_in = Ein_bitmap32[y_32][31-x_32];
                                            end
                                            [344:375]: begin        // D
                                                x_32 = x_pixel - (344);
                                                font_out = Dout_bitmap32[y_32][31-x_32];
                                                Y_in = Din_bitmap32[y_32][31-x_32];
                                            end
                                        endcase
                                end //red
                                2'd2: begin     //YELLOW
                                        case (x_pixel) inside
                                            [264:295]: begin        // Y
                                                x_32 = x_pixel - (264);
                                                font_out = Yout_bitmap32[y_32][31-x_32];
                                                G_in = Yin_bitmap32[y_32][31-x_32];
                                            end
                                            [304:335]: begin        // E
                                                x_32 = x_pixel - (304);
                                                font_out = Eout_bitmap32[y_32][31-x_32];
                                                G_in = Ein_bitmap32[y_32][31-x_32];
                                            end
                                            [344:375]: begin        // L
                                                x_32 = x_pixel - (344);
                                                font_out = Lout_bitmap32[y_32][31-x_32];
                                                G_in = Lin_bitmap32[y_32][31-x_32];
                                            end
                                        endcase
                                end
                                2'd3: begin     //YELLOW
                                        case (x_pixel) inside
                                            [264:295]: begin        // B
                                                x_32 = x_pixel - (264);
                                                font_out = Bout_bitmap32[y_32][31-x_32];
                                                R_in = Bin_bitmap32[y_32][31-x_32];
                                            end
                                            [304:335]: begin        // L
                                                x_32 = x_pixel - (304);
                                                font_out = Lout_bitmap32[y_32][31-x_32];
                                                R_in = Lin_bitmap32[y_32][31-x_32];
                                            end
                                            [344:375]: begin        // U
                                                x_32 = x_pixel - (344);
                                                font_out = Uout_bitmap32[y_32][31-x_32];
                                                R_in = Uin_bitmap32[y_32][31-x_32];
                                            end
                                        endcase
                                end //blue
                            endcase
                        end
                        [450:570]: begin
                            case (question[5:4])
                                2'd0: {red_port, green_port, blue_port} = {4'h0, 4'h0, 4'h0}; //black 0 들어오면 검정색
                                2'd1: begin     // BLUE
                                        case (x_pixel) inside
                                            [454:485]: begin        // R
                                                x_32 = x_pixel - (454);
                                                font_out = Rout_bitmap32[y_32][31-x_32];
                                                P_in = Rin_bitmap32[y_32][31-x_32];
                                            end
                                            [494:525]: begin        // E
                                                x_32 = x_pixel - (494);
                                                font_out = Eout_bitmap32[y_32][31-x_32];
                                                P_in = Ein_bitmap32[y_32][31-x_32];
                                            end
                                            [534:565]: begin        // D
                                                x_32 = x_pixel - (534);
                                                font_out = Dout_bitmap32[y_32][31-x_32];
                                                P_in = Din_bitmap32[y_32][31-x_32];
                                            end
                                        endcase
                                end //reR
                                2'd2: begin     // BLUE
                                        case (x_pixel) inside
                                            [454:485]: begin        // Y
                                                x_32 = x_pixel - (454);
                                                font_out = Yout_bitmap32[y_32][31-x_32];
                                                B_in = Yin_bitmap32[y_32][31-x_32];
                                            end
                                            [494:525]: begin        // E
                                                x_32 = x_pixel - (494);
                                                font_out = Eout_bitmap32[y_32][31-x_32];
                                                B_in = Ein_bitmap32[y_32][31-x_32];
                                            end
                                            [534:565]: begin        // L
                                                x_32 = x_pixel - (534);
                                                font_out = Lout_bitmap32[y_32][31-x_32];
                                                B_in = Lin_bitmap32[y_32][31-x_32];
                                            end
                                        endcase
                                end //yellow
                                2'd3: begin     // BLUE
                                        case (x_pixel) inside
                                            [454:485]: begin        // B
                                                x_32 = x_pixel - (454);
                                                font_out = Bout_bitmap32[y_32][31-x_32];
                                                G_in = Bin_bitmap32[y_32][31-x_32];
                                            end
                                            [494:525]: begin        // L
                                                x_32 = x_pixel - (494);
                                                font_out = Lout_bitmap32[y_32][31-x_32];
                                                G_in = Lin_bitmap32[y_32][31-x_32];
                                            end
                                            [534:565]: begin        // U
                                                x_32 = x_pixel - (534);
                                                font_out = Uout_bitmap32[y_32][31-x_32];
                                                G_in = Uin_bitmap32[y_32][31-x_32];
                                            end
                                        endcase
                                end
                            endcase
                        end
                        default: {red_port, green_port, blue_port} = {cam_r, cam_g, cam_b};
                        endcase 
                    end 
                 
                


                // 정답 제출할 영역 표시 (y= 280~400, x= 70 ~ 190), (y= 280~400, x= 260 ~ 380) , (y= 280~400, x= 450 ~ 570)
                else if (((x_pixel < 190 && x_pixel >= 70) && (y_pixel == 280 || y_pixel == 400)) ||
                        ((x_pixel == 190 || x_pixel == 70) && (y_pixel >= 280 && y_pixel < 400))) begin
                    red_port   = 4'h0;  
                    green_port = 4'h0;  
                    blue_port  = 4'h0;  // -> black 
                end else if (((x_pixel < 380 && x_pixel >= 260) && (y_pixel == 280 || y_pixel == 400)) ||
                            ((x_pixel == 380 || x_pixel == 260) && (y_pixel >= 280 && y_pixel < 400))) begin
                    red_port   = 4'h0;  
                    green_port = 4'h0;  
                    blue_port  = 4'h0;  // -> black  
                end else if (((x_pixel < 570 && x_pixel >= 450) && (y_pixel == 280 || y_pixel == 400)) ||
                            ((x_pixel == 570 || x_pixel == 450) && (y_pixel >= 280 && y_pixel < 400))) begin
                    red_port   = 4'h0;  
                    green_port = 4'h0;  
                    blue_port  = 4'h0;  // -> black  
                end 



                // LEVEL 3 표시 (y= 28~60, x= 210 ~ 436) 
                else if (y_pixel >= 28 && y_pixel < 60) begin
                    y_32 = y_pixel - 28;
                    case (x_pixel) inside
                        [210:241]: begin        // L
                            x_32 = x_pixel - (210);
                            font_out = Lout_bitmap32[y_32][31-x_32];
                            font_in = Lin_bitmap32[y_32][31-x_32];
                        end
                        [243:274]: begin        // E
                            x_32 = x_pixel - (243);
                            font_out = Eout_bitmap32[y_32][31-x_32];
                            font_in = Ein_bitmap32[y_32][31-x_32];
                        end
                        [276:307]: begin        // V
                            x_32 = x_pixel - (276);
                            font_out = Vout_bitmap32[y_32][31-x_32];
                            font_in = Vin_bitmap32[y_32][31-x_32];
                        end
                        [309:340]: begin        // E
                            x_32 = x_pixel - (309);
                            font_out = Eout_bitmap32[y_32][31-x_32];
                            font_in = Ein_bitmap32[y_32][31-x_32];
                        end
                        [342:373]: begin        // L
                            x_32 = x_pixel - (342);
                            font_out = Lout_bitmap32[y_32][31-x_32];
                            font_in = Lin_bitmap32[y_32][31-x_32];
                        end
                        [405:436]: begin        // 3
                            x_32 = x_pixel - (405);
                            font_out = threeout_bitmap32[y_32][31-x_32];
                            font_in = threein_bitmap32[y_32][31-x_32];
                        end
                        [440:471]: begin        // -
                            x_32 = x_pixel - (440);
                            font_out = dashout_bitmap32[y_32][31-x_32];
                            font_in = dashin_bitmap32[y_32][31-x_32];
                        end
                        [475:506]: begin        // 2
                            x_32 = x_pixel - (475);
                            font_out = twoout_bitmap32[y_32][31-x_32];
                            font_in = twoin_bitmap32[y_32][31-x_32];
                        end
                        [550:581]: begin       // countdown (y= 28~60, x=500~532 )
                        if (q_display_done) begin
                            x_32 = x_pixel - (550);
                            case (countdown)
                            4'd0: begin
                                font_out = zeroout_bitmap32[y_32][31-x_32];
                                countcolor_in = zeroin_bitmap32[y_32][31-x_32];
                            end 
                            4'd1: begin
                                font_out = oneout_bitmap32[y_32][31-x_32];
                                countcolor_in = onein_bitmap32[y_32][31-x_32];
                            end 
                            4'd2: begin
                                font_out = twoout_bitmap32[y_32][31-x_32];
                                countcolor_in = twoin_bitmap32[y_32][31-x_32];
                            end 
                            4'd3: begin
                                font_out = threeout_bitmap32[y_32][31-x_32];
                                countcolor_in = threein_bitmap32[y_32][31-x_32];
                            end 
                            4'd4: begin
                                font_out = fourout_bitmap32[y_32][31-x_32];
                                countcolor_in = fourin_bitmap32[y_32][31-x_32];
                            end 
                            4'd5: begin
                                font_out = fiveout_bitmap32[y_32][31-x_32];
                                countcolor_in = fivein_bitmap32[y_32][31-x_32];
                            end 
                            4'd6: begin
                                font_out = sixout_bitmap32[y_32][31-x_32];
                                countcolor_in = sixin_bitmap32[y_32][31-x_32];
                            end 
                            4'd7: begin
                                font_out = sevenout_bitmap32[y_32][31-x_32];
                                countcolor_in = sevenin_bitmap32[y_32][31-x_32];
                            end 
                            4'd8: begin
                                font_out = eightout_bitmap32[y_32][31-x_32];
                                countcolor_in = eightin_bitmap32[y_32][31-x_32];
                            end 
                            4'd9: begin
                                font_out = nineout_bitmap32[y_32][31-x_32];
                                countcolor_in = ninein_bitmap32[y_32][31-x_32];
                            end 
                            endcase
                        end
                        end
                    endcase
                end
                

                // 카운트 다운용 카운터 
                if (clk_counter == 25_000_000 - 1) begin
                    clk_counter_next = 0;  // 카운터 초기화
                    if (countdown > 0) begin
                        countdown_next = countdown - 1;  // 카운트다운 감소
                    end else begin
                        countdown_next = 0;  // 카운트다운이 0이 되면 유지
                    end
                end else begin
                    clk_counter_next = clk_counter + 1;  // 카운터 증가
                end

                if (countdown == 0) begin
                    countdown_done_next = 1;  // 카운트다운 완료 신호
                    q_display_done_next = 0;
                    // win 
                    state_next = WIN_LOSE;
                end 
            end

            LEVEL3_3: // Blink + 글자 4개 (글자와 색깔 다르게)
            begin
                // blink counter
                led_next = 4'b0100;
                if (clk_counter_blink == 2_500_000 - 1) begin
                    clk_counter_blink_next = 0;  // 카운터 초기화
                    if (blink_count == 49) begin
                        blink_count_next = 0;
                    end else begin
                        blink_count_next = blink_count + 1;
                    end
                end else begin
                    clk_counter_blink_next = clk_counter_blink + 1;  // 카운터 증가
                end



                 // 게임 색깔 표시 (4개) (y= 80~200, x= 32 ~ 152) , (y= 80~200, x= 184 ~ 304) , (y= 80~200, x= 336 ~ 456) , (y= 80~200, x= 488 ~ 608) 
                if (y_pixel >= 124 && y_pixel < 156) begin
                        y_32 = y_pixel - 124;
                        q_display_done_next = 1;
                        case (x_pixel) inside
                        [0:159]:begin
                            case (question[1:0])
                                2'd0: {red_port, green_port, blue_port} = {4'h0, 4'h0, 4'h0}; //black 0 들어오면 검정색
                                2'd1: begin     //RED
                                        case (x_pixel) inside
                                            [24:55]: begin        // R
                                                x_32 = x_pixel - (24);
                                                font_out = Rout_bitmap32[y_32][31-x_32];
                                                B_in = Rin_bitmap32[y_32][31-x_32];
                                            end
                                            [64:95]: begin        // E
                                                x_32 = x_pixel - (64);
                                                font_out = Eout_bitmap32[y_32][31-x_32];
                                                B_in = Ein_bitmap32[y_32][31-x_32];
                                            end
                                            [104:135]: begin        // D
                                                x_32 = x_pixel - (104);
                                                font_out = Dout_bitmap32[y_32][31-x_32];
                                                B_in = Din_bitmap32[y_32][31-x_32];
                                            end
                                        endcase
                                end
                                2'd2: case (x_pixel) inside
                                            [24:55]: begin        // Y
                                                x_32 = x_pixel - (24);
                                                font_out = Yout_bitmap32[y_32][31-x_32];
                                                G_in = Yin_bitmap32[y_32][31-x_32];
                                            end
                                            [64:95]: begin        // E
                                                x_32 = x_pixel - (64);
                                                font_out = Eout_bitmap32[y_32][31-x_32];
                                                G_in = Ein_bitmap32[y_32][31-x_32];
                                            end
                                            [104:135]: begin      // L
                                                x_32 = x_pixel - (104);
                                                font_out = Lout_bitmap32[y_32][31-x_32];
                                                G_in = Lin_bitmap32[y_32][31-x_32];
                                            end
                                        endcase //yellow
                                2'd3: case (x_pixel) inside
                                            [24:55]: begin        // B
                                                x_32 = x_pixel - (24);
                                                font_out = Bout_bitmap32[y_32][31-x_32];
                                                Y_in = Bin_bitmap32[y_32][31-x_32];
                                            end
                                            [64:95]: begin        // L
                                                x_32 = x_pixel - (64);
                                                font_out = Lout_bitmap32[y_32][31-x_32];
                                                Y_in = Lin_bitmap32[y_32][31-x_32];
                                            end
                                            [104:135]: begin      // U
                                                x_32 = x_pixel - (104);
                                                font_out = Uout_bitmap32[y_32][31-x_32];
                                                Y_in = Uin_bitmap32[y_32][31-x_32];
                                            end
                                        endcase //blue
                            endcase
                        end
                        [160:319]: begin
                            case (question[3:2])
                                2'd0: {red_port, green_port, blue_port} = {4'h0, 4'h0, 4'h0}; //black 0 들어오면 검정색
                                2'd1: begin     //YELLOW
                                        case (x_pixel) inside
                                            [184:215]: begin        // R
                                                x_32 = x_pixel - (184);
                                                font_out = Rout_bitmap32[y_32][31-x_32];
                                                Y_in = Rin_bitmap32[y_32][31-x_32];
                                            end
                                            [224:255]: begin        // E
                                                x_32 = x_pixel - (224);
                                                font_out = Eout_bitmap32[y_32][31-x_32];
                                                Y_in = Ein_bitmap32[y_32][31-x_32];
                                            end
                                            [264:295]: begin        // D
                                                x_32 = x_pixel - (264);
                                                font_out = Dout_bitmap32[y_32][31-x_32];
                                                Y_in = Din_bitmap32[y_32][31-x_32];
                                            end
                                        endcase
                                end //red
                                2'd2: begin     //YELLOW
                                        case (x_pixel) inside
                                            [184:215]: begin        // Y
                                                x_32 = x_pixel - (184);
                                                font_out = Yout_bitmap32[y_32][31-x_32];
                                                R_in = Yin_bitmap32[y_32][31-x_32];
                                            end
                                            [224:255]: begin        // E
                                                x_32 = x_pixel - (224);
                                                font_out = Eout_bitmap32[y_32][31-x_32];
                                                R_in = Ein_bitmap32[y_32][31-x_32];
                                            end
                                            [264:295]: begin        // L
                                                x_32 = x_pixel - (264);
                                                font_out = Lout_bitmap32[y_32][31-x_32];
                                                R_in = Lin_bitmap32[y_32][31-x_32];
                                            end
                                        endcase
                                end
                                2'd3: begin     //YELLOW
                                        case (x_pixel) inside
                                            [184:215]: begin        // B
                                                x_32 = x_pixel - (184);
                                                font_out = Bout_bitmap32[y_32][31-x_32];
                                                P_in = Bin_bitmap32[y_32][31-x_32];
                                            end
                                            [224:255]: begin        // L
                                                x_32 = x_pixel - (224);
                                                font_out = Lout_bitmap32[y_32][31-x_32];
                                                P_in = Lin_bitmap32[y_32][31-x_32];
                                            end
                                            [264:295]: begin        // U
                                                x_32 = x_pixel - (264);
                                                font_out = Uout_bitmap32[y_32][31-x_32];
                                                P_in = Uin_bitmap32[y_32][31-x_32];
                                            end
                                        endcase
                                end //blue
                            endcase
                        end
                        [320:479]: begin
                            case (question[5:4])
                                2'd0: {red_port, green_port, blue_port} = {4'h0, 4'h0, 4'h0}; //black 0 들어오면 검정색
                                2'd1: begin     // BLU
                                        case (x_pixel) inside
                                            [344:375]: begin        // R
                                                x_32 = x_pixel - (344);
                                                font_out = Rout_bitmap32[y_32][31-x_32];
                                                P_in = Rin_bitmap32[y_32][31-x_32];
                                            end
                                            [384:415]: begin        // E
                                                x_32 = x_pixel - (384);
                                                font_out = Eout_bitmap32[y_32][31-x_32];
                                                P_in = Ein_bitmap32[y_32][31-x_32];
                                            end
                                            [424:455]: begin        // D
                                                x_32 = x_pixel - (424);
                                                font_out = Dout_bitmap32[y_32][31-x_32];
                                                P_in = Din_bitmap32[y_32][31-x_32];
                                            end
                                        endcase
                                end //red
                                2'd2: begin     // BLUE
                                        case (x_pixel) inside
                                            [344:375]: begin        // Y
                                                x_32 = x_pixel - (344);
                                                font_out = Yout_bitmap32[y_32][31-x_32];
                                                B_in = Yin_bitmap32[y_32][31-x_32];
                                            end
                                            [384:415]: begin        // E
                                                x_32 = x_pixel - (384);
                                                font_out = Eout_bitmap32[y_32][31-x_32];
                                                B_in = Ein_bitmap32[y_32][31-x_32];
                                            end
                                            [424:455]: begin        // L
                                                x_32 = x_pixel - (424);
                                                font_out = Lout_bitmap32[y_32][31-x_32];
                                                B_in = Lin_bitmap32[y_32][31-x_32];
                                            end
                                        endcase
                                end //yellow
                                2'd3: begin     // BLUE
                                        case (x_pixel) inside
                                            [344:375]: begin        // B
                                                x_32 = x_pixel - (344);
                                                font_out = Bout_bitmap32[y_32][31-x_32];
                                                G_in = Bin_bitmap32[y_32][31-x_32];
                                            end
                                            [384:415]: begin        // L
                                                x_32 = x_pixel - (384);
                                                font_out = Lout_bitmap32[y_32][31-x_32];
                                                G_in = Lin_bitmap32[y_32][31-x_32];
                                            end
                                            [424:455]: begin        // U
                                                x_32 = x_pixel - (424);
                                                font_out = Uout_bitmap32[y_32][31-x_32];
                                                G_in = Uin_bitmap32[y_32][31-x_32];
                                            end
                                        endcase
                                end
                            endcase
                        end
                        [480:639]:begin
                            case (question[7:6])
                                2'd0: {red_port, green_port, blue_port} = {4'h0, 4'h0, 4'h0}; //black 0 들어오면 검정색
                                2'd1: begin     //RED
                                        case (x_pixel) inside
                                            [504:535]: begin        // R
                                                x_32 = x_pixel - (504);
                                                font_out = Rout_bitmap32[y_32][31-x_32];
                                                G_in = Rin_bitmap32[y_32][31-x_32];
                                            end
                                            [544:575]: begin        // E
                                                x_32 = x_pixel - (544);
                                                font_out = Eout_bitmap32[y_32][31-x_32];
                                                G_in = Ein_bitmap32[y_32][31-x_32];
                                            end
                                            [584:615]: begin        // D
                                                x_32 = x_pixel - (584);
                                                font_out = Dout_bitmap32[y_32][31-x_32];
                                                G_in = Din_bitmap32[y_32][31-x_32];
                                            end
                                        endcase
                                end
                                2'd2: begin     //RED
                                        case (x_pixel) inside
                                            [504:535]: begin        // Y
                                                x_32 = x_pixel - (504);
                                                font_out = Yout_bitmap32[y_32][31-x_32];
                                                P_in = Yin_bitmap32[y_32][31-x_32];
                                            end
                                            [544:575]: begin        // E
                                                x_32 = x_pixel - (544);
                                                font_out = Eout_bitmap32[y_32][31-x_32];
                                                P_in = Ein_bitmap32[y_32][31-x_32];
                                            end
                                            [584:615]: begin        // L
                                                x_32 = x_pixel - (584);
                                                font_out = Lout_bitmap32[y_32][31-x_32];
                                                P_in = Lin_bitmap32[y_32][31-x_32];
                                            end
                                        endcase
                                end //yellow
                                2'd3: begin     //RED
                                        case (x_pixel) inside
                                            [504:535]: begin        // B
                                                x_32 = x_pixel - (504);
                                                font_out = Bout_bitmap32[y_32][31-x_32];
                                                R_in = Bin_bitmap32[y_32][31-x_32];
                                            end
                                            [544:575]: begin        // L
                                                x_32 = x_pixel - (544);
                                                font_out = Lout_bitmap32[y_32][31-x_32];
                                                R_in = Lin_bitmap32[y_32][31-x_32];
                                            end
                                            [584:615]: begin        // U
                                                x_32 = x_pixel - (584);
                                                font_out = Uout_bitmap32[y_32][31-x_32];
                                                R_in = Uin_bitmap32[y_32][31-x_32];
                                            end
                                        endcase
                                end //blue
                            endcase     
                        end
                        default: {red_port, green_port, blue_port} = {cam_r, cam_g, cam_b};
                        endcase 
                    end 
                 
                


                // 정답 제출할 영역 표시 (y= 280~400, x= 32 ~ 152), (y= 280~400, x= 184 ~ 304) , (y= 280~400, x= 336 ~ 456)  , (y= 280~400, x= 488 ~ 608)  
                else if (((x_pixel < 152 && x_pixel >= 32) && (y_pixel == 280 || y_pixel == 400)) ||
                        ((x_pixel == 152 || x_pixel == 32) && (y_pixel >= 280 && y_pixel < 400))) begin
                    red_port   = 4'h0;  
                    green_port = 4'h0;  
                    blue_port  = 4'h0;  // -> black 
                end else if (((x_pixel < 304 && x_pixel >= 184) && (y_pixel == 280 || y_pixel == 400)) ||
                            ((x_pixel == 304 || x_pixel == 184) && (y_pixel >= 280 && y_pixel < 400))) begin
                    red_port   = 4'h0;  
                    green_port = 4'h0;  
                    blue_port  = 4'h0;  // -> black  
                end else if (((x_pixel < 456 && x_pixel >= 336) && (y_pixel == 280 || y_pixel == 400)) ||
                            ((x_pixel == 456 || x_pixel == 336) && (y_pixel >= 280 && y_pixel < 400))) begin
                    red_port   = 4'h0;  
                    green_port = 4'h0;  
                    blue_port  = 4'h0;  // -> black  
                end else if (((x_pixel < 608 && x_pixel >= 488) && (y_pixel == 280 || y_pixel == 400)) ||
                            ((x_pixel == 608 || x_pixel == 488) && (y_pixel >= 280 && y_pixel < 400))) begin
                    red_port   = 4'h0;  
                    green_port = 4'h0;  
                    blue_port  = 4'h0;  // -> black  
                end 



                // LEVEL 3 표시 (y= 28~60, x= 210 ~ 436) 
                else if (y_pixel >= 28 && y_pixel < 60) begin
                    y_32 = y_pixel - 28;
                    case (x_pixel) inside
                        [210:241]: begin        // L
                            x_32 = x_pixel - (210);
                            font_out = Lout_bitmap32[y_32][31-x_32];
                            font_in = Lin_bitmap32[y_32][31-x_32];
                        end
                        [243:274]: begin        // E
                            x_32 = x_pixel - (243);
                            font_out = Eout_bitmap32[y_32][31-x_32];
                            font_in = Ein_bitmap32[y_32][31-x_32];
                        end
                        [276:307]: begin        // V
                            x_32 = x_pixel - (276);
                            font_out = Vout_bitmap32[y_32][31-x_32];
                            font_in = Vin_bitmap32[y_32][31-x_32];
                        end
                        [309:340]: begin        // E
                            x_32 = x_pixel - (309);
                            font_out = Eout_bitmap32[y_32][31-x_32];
                            font_in = Ein_bitmap32[y_32][31-x_32];
                        end
                        [342:373]: begin        // L
                            x_32 = x_pixel - (342);
                            font_out = Lout_bitmap32[y_32][31-x_32];
                            font_in = Lin_bitmap32[y_32][31-x_32];
                        end
                        [405:436]: begin        // 3
                            x_32 = x_pixel - (405);
                            font_out = threeout_bitmap32[y_32][31-x_32];
                            font_in = threein_bitmap32[y_32][31-x_32];
                        end
                        [440:471]: begin        // -
                            x_32 = x_pixel - (440);
                            font_out = dashout_bitmap32[y_32][31-x_32];
                            font_in = dashin_bitmap32[y_32][31-x_32];
                        end
                        [475:506]: begin        // 3
                            x_32 = x_pixel - (475);
                            font_out = threeout_bitmap32[y_32][31-x_32];
                            font_in = threein_bitmap32[y_32][31-x_32];
                        end
                        [550:581]: begin       // countdown (y= 28~60, x=500~532 )
                        if (q_display_done) begin
                            x_32 = x_pixel - (550);
                            case (countdown)
                            4'd0: begin
                                font_out = zeroout_bitmap32[y_32][31-x_32];
                                countcolor_in = zeroin_bitmap32[y_32][31-x_32];
                            end 
                            4'd1: begin
                                font_out = oneout_bitmap32[y_32][31-x_32];
                                countcolor_in = onein_bitmap32[y_32][31-x_32];
                            end 
                            4'd2: begin
                                font_out = twoout_bitmap32[y_32][31-x_32];
                                countcolor_in = twoin_bitmap32[y_32][31-x_32];
                            end 
                            4'd3: begin
                                font_out = threeout_bitmap32[y_32][31-x_32];
                                countcolor_in = threein_bitmap32[y_32][31-x_32];
                            end 
                            4'd4: begin
                                font_out = fourout_bitmap32[y_32][31-x_32];
                                countcolor_in = fourin_bitmap32[y_32][31-x_32];
                            end 
                            4'd5: begin
                                font_out = fiveout_bitmap32[y_32][31-x_32];
                                countcolor_in = fivein_bitmap32[y_32][31-x_32];
                            end 
                            4'd6: begin
                                font_out = sixout_bitmap32[y_32][31-x_32];
                                countcolor_in = sixin_bitmap32[y_32][31-x_32];
                            end 
                            4'd7: begin
                                font_out = sevenout_bitmap32[y_32][31-x_32];
                                countcolor_in = sevenin_bitmap32[y_32][31-x_32];
                            end 
                            4'd8: begin
                                font_out = eightout_bitmap32[y_32][31-x_32];
                                countcolor_in = eightin_bitmap32[y_32][31-x_32];
                            end 
                            4'd9: begin
                                font_out = nineout_bitmap32[y_32][31-x_32];
                                countcolor_in = ninein_bitmap32[y_32][31-x_32];
                            end 
                            endcase
                        end
                        end
                    endcase
                end
                

                // 카운트 다운용 카운터 
                if (clk_counter == 25_000_000 - 1) begin
                    clk_counter_next = 0;  // 카운터 초기화
                    if (countdown > 0) begin
                        countdown_next = countdown - 1;  // 카운트다운 감소
                    end else begin
                        countdown_next = 0;  // 카운트다운이 0이 되면 유지
                    end
                end else begin
                    clk_counter_next = clk_counter + 1;  // 카운터 증가
                end

                if (countdown == 0) begin
                    countdown_done_next = 1;  // 카운트다운 완료 신호
                    q_display_done_next = 0;
                    // win 
                    state_next = WIN_LOSE;
                end 
            end

  




        /************************************WIN_LOSE******************************************/
        /************************************WIN_LOSE******************************************/
        /************************************WIN_LOSE******************************************/
        /************************************WIN_LOSE******************************************/
        /************************************WIN_LOSE******************************************/
        /************************************WIN_LOSE******************************************/
        /************************************WIN_LOSE******************************************/
        /************************************WIN_LOSE******************************************/
        /************************************WIN_LOSE******************************************/
        /************************************WIN_LOSE******************************************/
        WIN_LOSE : begin
            countdown_done_next = 0;
            led_next = 4'b1111;
            temp_y_coordinate_next = WL_DISPLAY_Y1;
            if (comparison_done) begin
                give_comparison_done_next = 1;
                if (win_lose == 2'b01) begin 
                    // 받았다고 보내기
                    state_next = WIN_DSIPLAY;
                    countdown_done_next = 0;
                    score_next = score + 1;
                    
                    
                // lose 표시
                end else if (win_lose == 2'b10) begin  
                    state_next = LOSE_DSIPLAY;
                    countdown_done_next = 0;
                    
                
                end else begin
                    countdown_done_next = 0;
                end
            end else begin
                    countdown_done_next = 0;
            end
        end


        /************************************WIN_DISPLAY******************************************/
        /************************************WIN_DISPLAY******************************************/
        /************************************WIN_DISPLAY******************************************/
        /************************************WIN_DISPLAY******************************************/
        /************************************WIN_DISPLAY******************************************/
        /************************************WIN_DISPLAY******************************************/
        /************************************WIN_DISPLAY******************************************/
        /************************************WIN_DISPLAY******************************************/
        /************************************WIN_DISPLAY******************************************/
        /************************************WIN_DISPLAY******************************************/
        WIN_DSIPLAY : 
        
        begin
            give_comparison_done_next = 0;

            if ((y_pixel >= WL_DISPLAY_Y1) && (y_pixel < (WL_DISPLAY_Y1 + WIDTH64))) begin
                    y_64 = y_pixel - WL_DISPLAY_Y1;
                    //win display

                    case (x_pixel) inside
                        [W_X_COORDINATE : W_X_COORDINATE + WIDTH64 - 1]: begin
                            x_64 = x_pixel - W_X_COORDINATE;
                            w_out = Wout_bitmap[y_64][63-x_64];
                            w_mid = Wmid_bitmap[y_64][63-x_64];
                            w_in = Win_bitmap[y_64][63-x_64];
                        end
                        [(W_X_COORDINATE + WIDTH64 + LETTER_INTERVAL) : (W_X_COORDINATE + WIDTH64 + WIDTH32 + LETTER_INTERVAL) - 1]: begin
                            x_32 = x_pixel - (W_X_COORDINATE + WIDTH64 + LETTER_INTERVAL);
                            w_out = i1_bitmap[y_64][31-x_32];
                            w_mid = i2_bitmap[y_64][31-x_32];
                            w_in = i3_bitmap[y_64][31-x_32];
                        end
                        [(W_X_COORDINATE + WIDTH64 + WIDTH32 + 2*LETTER_INTERVAL) : (W_X_COORDINATE + 2*WIDTH64 + WIDTH32 + 2*LETTER_INTERVAL) - 1]: begin
                            x_64 = x_pixel - (W_X_COORDINATE + WIDTH64 + WIDTH32 + 2*LETTER_INTERVAL);
                            w_out = n1_bitmap[y_64][63-x_64];
                            w_mid = n2_bitmap[y_64][63-x_64];
                            w_in = n3_bitmap[y_64][63-x_64];
                        end
                        [(W_X_COORDINATE + 2*WIDTH64 + WIDTH32 + 3*LETTER_INTERVAL) : (W_X_COORDINATE + 2*WIDTH64 + 2*WIDTH32 + 3*LETTER_INTERVAL) - 1]: begin
                            x_32 = x_pixel - (W_X_COORDINATE + 2*WIDTH64 + WIDTH32 + 3*LETTER_INTERVAL);
                            w_out = ex1_bitmap[y_64][31-x_32];
                            w_mid = ex2_bitmap[y_64][31-x_32];
                            w_in = ex3_bitmap[y_64][31-x_32];
                        end
                        [(W_X_COORDINATE + 2*WIDTH64 + 2*WIDTH32 + 4*LETTER_INTERVAL) : (W_X_COORDINATE + 2*WIDTH64 + 3*WIDTH32 + 4*LETTER_INTERVAL) - 1]: begin
                            x_32 = x_pixel - (W_X_COORDINATE + 2*WIDTH64 + 2*WIDTH32 + 4*LETTER_INTERVAL);
                            w_out = ex1_bitmap[y_64][31-x_32];
                            w_mid = ex2_bitmap[y_64][31-x_32];
                            w_in = ex3_bitmap[y_64][31-x_32];
                        end
                    endcase

                    if ( (y_pixel >= (WL_DISPLAY_Y1 + 16)) && (y_pixel < (WL_DISPLAY_Y1 + 48))) begin
                        y_32 = y_pixel - (WL_DISPLAY_Y1 + 16);
                        case (x_pixel) inside
                            [(SCORE_X_COORDINATE):(SCORE_X_COORDINATE + WIDTH32) -1 ]: begin
                            x_32 = x_pixel - (SCORE_X_COORDINATE);
                            case (score / 10)
                                4'd0: begin
                                    font_out = zeroout_bitmap32[y_32][31-x_32];
                                    font_in  = zeroin_bitmap32[y_32][31-x_32];                    
                                end

                                4'd1: begin
                                    font_out = oneout_bitmap32[y_32][31-x_32];
                                    font_in  = onein_bitmap32[y_32][31-x_32];                    
                                end

                                4'd2: begin
                                    font_out = twoout_bitmap32[y_32][31-x_32];
                                    font_in  = twoin_bitmap32[y_32][31-x_32];                    
                                end

                                4'd3: begin
                                    font_out = threeout_bitmap32[y_32][31-x_32];
                                    font_in  = threein_bitmap32[y_32][31-x_32];                    
                                end

                                4'd4: begin
                                    font_out = fourout_bitmap32[y_32][31-x_32];
                                    font_in  = fourin_bitmap32[y_32][31-x_32];                    
                                end

                                4'd5: begin
                                    font_out = fiveout_bitmap32[y_32][31-x_32];
                                    font_in  = fivein_bitmap32[y_32][31-x_32];                    
                                end

                                4'd6: begin
                                    font_out = sixout_bitmap32[y_32][31-x_32];
                                    font_in  = sixin_bitmap32[y_32][31-x_32];                    
                                end

                                4'd7: begin
                                    font_out = sevenout_bitmap32[y_32][31-x_32];
                                    font_in  = sevenin_bitmap32[y_32][31-x_32];                    
                                end

                                4'd8: begin
                                    font_out = eightout_bitmap32[y_32][31-x_32];
                                    font_in  = eightin_bitmap32[y_32][31-x_32];                    
                                end

                                4'd9: begin
                                    font_out = nineout_bitmap32[y_32][31-x_32];
                                    font_in  = ninein_bitmap32[y_32][31-x_32];                    
                                end

                                default: begin
                                    font_out = zeroout_bitmap32[y_32][31-x_32];
                                    font_in  = zeroin_bitmap32[y_32][31-x_32];                                        
                                end
                            endcase
                            end
                            [(SCORE_X_COORDINATE + WIDTH32 ):(SCORE_X_COORDINATE + 2*WIDTH32 )-1]: begin
                            x_32 = x_pixel - (SCORE_X_COORDINATE + WIDTH32 );
                            case (score % 10)
                                4'd0: begin
                                    font_out = zeroout_bitmap32[y_32][31-x_32];
                                    font_in  = zeroin_bitmap32[y_32][31-x_32];                    
                                end

                                4'd1: begin
                                    font_out = oneout_bitmap32[y_32][31-x_32];
                                    font_in  = onein_bitmap32[y_32][31-x_32];                    
                                end

                                4'd2: begin
                                    font_out = twoout_bitmap32[y_32][31-x_32];
                                    font_in  = twoin_bitmap32[y_32][31-x_32];                    
                                end

                                4'd3: begin
                                    font_out = threeout_bitmap32[y_32][31-x_32];
                                    font_in  = threein_bitmap32[y_32][31-x_32];                    
                                end

                                4'd4: begin
                                    font_out = fourout_bitmap32[y_32][31-x_32];
                                    font_in  = fourin_bitmap32[y_32][31-x_32];                    
                                end

                                4'd5: begin
                                    font_out = fiveout_bitmap32[y_32][31-x_32];
                                    font_in  = fivein_bitmap32[y_32][31-x_32];                    
                                end

                                4'd6: begin
                                    font_out = sixout_bitmap32[y_32][31-x_32];
                                    font_in  = sixin_bitmap32[y_32][31-x_32];                    
                                end

                                4'd7: begin
                                    font_out = sevenout_bitmap32[y_32][31-x_32];
                                    font_in  = sevenin_bitmap32[y_32][31-x_32];                    
                                end

                                4'd8: begin
                                    font_out = eightout_bitmap32[y_32][31-x_32];
                                    font_in  = eightin_bitmap32[y_32][31-x_32];                    
                                end

                                4'd9: begin
                                    font_out = nineout_bitmap32[y_32][31-x_32];
                                    font_in  = ninein_bitmap32[y_32][31-x_32];                    
                                end

                                default: begin
                                    font_out = zeroout_bitmap32[y_32][31-x_32];
                                    font_in  = zeroin_bitmap32[y_32][31-x_32];                                        
                                end
                            endcase     
                            end
                        endcase
                    end
                end 
                

                        if (clk_counter_delay == 25_000_000 - 1) begin
                            clk_counter_delay_next = 0;  // 카운터 초기화
                            if (delay_count == 10) begin
                                delay_count_next = 0;
                            end else begin
                                delay_count_next = delay_count + 1;
                            end
                        end else begin
                            clk_counter_delay_next = clk_counter_delay + 1;  // 카운터 증가
                        end

                        if (delay_count == 4) begin
                            game_done_next = 1;  // 게임 완료 신호 
                            delay_count_next = 0;
                            clk_counter_delay_next = 0;
                            frame_counter_next = 0;
                            frame_next = 0;
                            state_next = GAME_DONE;  // 다음 레벨로 이동
                        end         
            
                    end

        /************************************LOSE_DISPLAY******************************************/
        /************************************LOSE_DISPLAY******************************************/
        /************************************LOSE_DISPLAY******************************************/
        /************************************LOSE_DISPLAY******************************************/
        /************************************LOSE_DISPLAY******************************************/
        /************************************LOSE_DISPLAY******************************************/
        /************************************LOSE_DISPLAY******************************************/
        /************************************LOSE_DISPLAY******************************************/
        /************************************LOSE_DISPLAY******************************************/
        /************************************LOSE_DISPLAY******************************************/
        LOSE_DSIPLAY: 
        begin
            give_comparison_done_next = 0;
            //LOSE띄우기
             if ((y_pixel >= WL_DISPLAY_Y1) && (y_pixel < (WL_DISPLAY_Y1 + WIDTH64))) begin
                    y_64 = y_pixel - WL_DISPLAY_Y1;
                    
                    //win display

                    case (x_pixel) inside
                        [L_X_COORDINATE : (L_X_COORDINATE + WIDTH64) - 1]: begin
                             x_64 = x_pixel - L_X_COORDINATE;
                        L_mid = Lmid_bitmap[y_64][63 - x_64];
                        L_in  = Lin_bitmap[y_64][63 - x_64];
                        L_out = Lout_bitmap[y_64][63 - x_64];
                        end
                        [(L_X_COORDINATE + WIDTH64 + LETTER_INTERVAL) : (L_X_COORDINATE + 2*WIDTH64 + LETTER_INTERVAL) - 1]: begin
                            x_64 = x_pixel - (L_X_COORDINATE + WIDTH64 + LETTER_INTERVAL);
                        L_mid = Omid_bitmap[y_64][63 - x_64];
                        L_in  = Oin_bitmap[y_64][63 - x_64];
                        L_out = Oout_bitmap[y_64][63 - x_64];
                        end
                        [(L_X_COORDINATE + 2*WIDTH64 + 2*LETTER_INTERVAL) : (L_X_COORDINATE + 3*WIDTH64 + 2*LETTER_INTERVAL) - 1]: begin
                        x_64 = x_pixel - (L_X_COORDINATE + 2*WIDTH64 + 2*LETTER_INTERVAL);
                        L_mid = Smid_bitmap[y_64][63 - x_64];
                        L_in  = Sin_bitmap[y_64][63 - x_64];
                        L_out = Sout_bitmap[y_64][63 - x_64];
                        end
                        [(L_X_COORDINATE + 3*WIDTH64 + 3*LETTER_INTERVAL) : (L_X_COORDINATE + 4*WIDTH64 + 3*LETTER_INTERVAL) - 1]: begin
                         x_64 = x_pixel - (L_X_COORDINATE + 3*WIDTH64 + 3*LETTER_INTERVAL);
                        L_mid = Emid_bitmap[y_64][63 - x_64];
                        L_in  = Ein_bitmap[y_64][63 - x_64];
                        L_out = Eout_bitmap[y_64][63 - x_64];
                        end
                        [(L_X_COORDINATE + 4*WIDTH64 + 4*LETTER_INTERVAL) : (L_X_COORDINATE + 4*WIDTH64 + WIDTH32 + 4*LETTER_INTERVAL) - 1]: begin
                         x_32 = x_pixel - (L_X_COORDINATE + 4*WIDTH64 + 4*LETTER_INTERVAL);
                        L_out = ex1_bitmap[y_64][31-x_32];
                        L_mid = ex2_bitmap[y_64][31-x_32];
                        L_in = ex3_bitmap[y_64][31-x_32];
                        end
                        [(L_X_COORDINATE + 4*WIDTH64 + WIDTH32 + 5*LETTER_INTERVAL) : (L_X_COORDINATE + 4*WIDTH64 + 2*WIDTH32 + 5*LETTER_INTERVAL) - 1]: begin
                        x_32 = x_pixel - (L_X_COORDINATE + 4*WIDTH64 + WIDTH32 + 5*LETTER_INTERVAL);
                        L_out = ex1_bitmap[y_64][31-x_32];
                        L_mid = ex2_bitmap[y_64][31-x_32];
                        L_in = ex3_bitmap[y_64][31-x_32];
                        end
                    endcase

                    //score display
                if ( (y_pixel >= WL_DISPLAY_Y1 + 16) && (y_pixel < (WL_DISPLAY_Y1 + 48))) begin
                        y_32 = y_pixel - (WL_DISPLAY_Y1 + 16);
                        case (x_pixel) inside
                            [(SCORE_X_COORDINATE):(SCORE_X_COORDINATE + WIDTH32) -1 ]: begin
                            x_32 = x_pixel - (SCORE_X_COORDINATE);
                            case (score / 10)
                                4'd0: begin
                                    font_out = zeroout_bitmap32[y_32][31-x_32];
                                    font_in  = zeroin_bitmap32[y_32][31-x_32];                    
                                end

                                4'd1: begin
                                    font_out = oneout_bitmap32[y_32][31-x_32];
                                    font_in  = onein_bitmap32[y_32][31-x_32];                    
                                end

                                4'd2: begin
                                    font_out = twoout_bitmap32[y_32][31-x_32];
                                    font_in  = twoin_bitmap32[y_32][31-x_32];                    
                                end

                                4'd3: begin
                                    font_out = threeout_bitmap32[y_32][31-x_32];
                                    font_in  = threein_bitmap32[y_32][31-x_32];                    
                                end

                                4'd4: begin
                                    font_out = fourout_bitmap32[y_32][31-x_32];
                                    font_in  = fourin_bitmap32[y_32][31-x_32];                    
                                end

                                4'd5: begin
                                    font_out = fiveout_bitmap32[y_32][31-x_32];
                                    font_in  = fivein_bitmap32[y_32][31-x_32];                    
                                end

                                4'd6: begin
                                    font_out = sixout_bitmap32[y_32][31-x_32];
                                    font_in  = sixin_bitmap32[y_32][31-x_32];                    
                                end

                                4'd7: begin
                                    font_out = sevenout_bitmap32[y_32][31-x_32];
                                    font_in  = sevenin_bitmap32[y_32][31-x_32];                    
                                end

                                4'd8: begin
                                    font_out = eightout_bitmap32[y_32][31-x_32];
                                    font_in  = eightin_bitmap32[y_32][31-x_32];                    
                                end

                                4'd9: begin
                                    font_out = nineout_bitmap32[y_32][31-x_32];
                                    font_in  = ninein_bitmap32[y_32][31-x_32];                    
                                end

                                default: begin
                                    font_out = zeroout_bitmap32[y_32][31-x_32];
                                    font_in  = zeroin_bitmap32[y_32][31-x_32];                                        
                                end
                            endcase
                            end
                            [(SCORE_X_COORDINATE + WIDTH32 ):(SCORE_X_COORDINATE + 2*WIDTH32 )-1]: begin
                            x_32 = x_pixel - (SCORE_X_COORDINATE + WIDTH32 );
                            case (score % 10)
                                4'd0: begin
                                    font_out = zeroout_bitmap32[y_32][31-x_32];
                                    font_in  = zeroin_bitmap32[y_32][31-x_32];                    
                                end

                                4'd1: begin
                                    font_out = oneout_bitmap32[y_32][31-x_32];
                                    font_in  = onein_bitmap32[y_32][31-x_32];                    
                                end

                                4'd2: begin
                                    font_out = twoout_bitmap32[y_32][31-x_32];
                                    font_in  = twoin_bitmap32[y_32][31-x_32];                    
                                end

                                4'd3: begin
                                    font_out = threeout_bitmap32[y_32][31-x_32];
                                    font_in  = threein_bitmap32[y_32][31-x_32];                    
                                end

                                4'd4: begin
                                    font_out = fourout_bitmap32[y_32][31-x_32];
                                    font_in  = fourin_bitmap32[y_32][31-x_32];                    
                                end

                                4'd5: begin
                                    font_out = fiveout_bitmap32[y_32][31-x_32];
                                    font_in  = fivein_bitmap32[y_32][31-x_32];                    
                                end

                                4'd6: begin
                                    font_out = sixout_bitmap32[y_32][31-x_32];
                                    font_in  = sixin_bitmap32[y_32][31-x_32];                    
                                end

                                4'd7: begin
                                    font_out = sevenout_bitmap32[y_32][31-x_32];
                                    font_in  = sevenin_bitmap32[y_32][31-x_32];                    
                                end

                                4'd8: begin
                                    font_out = eightout_bitmap32[y_32][31-x_32];
                                    font_in  = eightin_bitmap32[y_32][31-x_32];                    
                                end

                                4'd9: begin
                                    font_out = nineout_bitmap32[y_32][31-x_32];
                                    font_in  = ninein_bitmap32[y_32][31-x_32];                    
                                end

                                default: begin
                                    font_out = zeroout_bitmap32[y_32][31-x_32];
                                    font_in  = zeroin_bitmap32[y_32][31-x_32];                                        
                                end
                            endcase     
                            end
                        endcase
                    end
                end
            
                if (clk_counter_delay == 25_000_000 - 1) begin
                    clk_counter_delay_next = 0;  // 카운터 초기화
                    if (delay_count == 10) begin
                        delay_count_next = 0;
                    end else begin
                        delay_count_next = delay_count + 1;
                    end
                end else begin
                    clk_counter_delay_next = clk_counter_delay + 1;  // 카운터 증가
                end

                if (delay_count == 4) begin
                    game_done_next = 1;  // 게임 완료 신호 
                    delay_count_next = 0;
                    clk_counter_delay_next = 0;
                    frame_counter_next = 0;
                    frame_next = 0;
                    state_next = GAME_DONE;  // 다음 레벨로 이동
                end 
                
            end



        /************************************GAME_DONE******************************************/
        /************************************GAME_DONE******************************************/
        /************************************GAME_DONE******************************************/
        /************************************GAME_DONE******************************************/
        /************************************GAME_DONE******************************************/
        /************************************GAME_DONE******************************************/
        /************************************GAME_DONE******************************************/
        /************************************GAME_DONE******************************************/
        /************************************GAME_DONE******************************************/
        /************************************GAME_DONE******************************************/
        /************************************GAME_DONE******************************************/
        /************************************GAME_DONE******************************************/
        /************************************GAME_DONE******************************************/


        GAME_DONE : 
            begin   
            // 이 상태에서 count_down이랑 blink count 초기화해줌
                if (give_done_ff2) begin 
                    blink_count_next = 0;
                    countdown_next = 5; 
                    state_next = HOLD;
                    game_done_next = 0;
                end 
            end

        HOLD : begin
            if(!give_done_ff2) begin
                if (end_reg) begin
                    end_next = 0;
                    countdown_next = 10;
                    state_next = END_DISPLAY;
                    game_done_next = 1;
                end else begin
                    state_next = SEL_LEVEL; 
                    game_done_next = 1;
                end
            end
        end
        
        SEL_LEVEL: // 레벨 받으면 각 레벨 상태로 이동 
             begin
                //lvl_count_next = lvl_count + 1;
                game_done_next = 1;
                led_next = 4'b0110;
                if (start_ff2) begin
                    case (lvl)
                        2'b00: state_next = LEVEL0;
                        2'b01: begin
                        if (lvl_count == 0) begin
                            state_next = LEVEL1_1;
                        end else if (lvl_count == 1) begin
                            state_next = LEVEL2_1;
                        end else if (lvl_count == 2) begin
                            state_next = LEVEL3_1;
                        end
                        end 
                        2'b10: begin
                        if (lvl_count == 0) begin
                            state_next = LEVEL1_2;
                        end else if (lvl_count == 1) begin
                            state_next = LEVEL2_2;
                        end else if (lvl_count == 2) begin
                            state_next = LEVEL3_2;
                        end
                        end 
                        2'b11:begin
                        if (lvl_count == 0) begin
                            lvl_count_next = lvl_count + 1;
                            state_next = LEVEL1_3;
                        end else if (lvl_count == 1) begin
                            lvl_count_next = lvl_count + 1;
                            state_next = LEVEL2_3;
                        end else if (lvl_count == 2) begin
                            lvl_count_next = 0;
                            state_next = LEVEL3_3;
                            end_next = 1;
                        end
                        end 
                    endcase
                end
            end

         END_DISPLAY :
            begin
                lvl_count_next = 0;     // 레벨 카운터 초기화
                game_done_next = 1;

                // THE END 표시
                if (y_pixel >= 80 && y_pixel < 112) begin
                    y_32 = y_pixel - 80;
                    case (x_pixel) inside
                        [204:235]: begin        // T
                            x_32 = x_pixel - (204);
                            font_out = Tout_bitmap32[y_32][31-x_32];
                            font_in = Tin_bitmap32[y_32][31-x_32];
                                            end
                        [238:269]: begin        // H
                            x_32 = x_pixel - (238);
                            font_out = Hout_bitmap32[y_32][31-x_32];
                            font_in = Hin_bitmap32[y_32][31-x_32];
                        end
                        [272:303]: begin        // E
                            x_32 = x_pixel - (272);
                            font_out = Eout_bitmap32[y_32][31-x_32];
                            font_in = Ein_bitmap32[y_32][31-x_32];
                        end
                        //space
                        [334:365]: begin        // E
                            x_32 = x_pixel - (334);
                            font_out = Eout_bitmap32[y_32][31-x_32];
                            font_in = Ein_bitmap32[y_32][31-x_32];
                                            end
                        [368:399]: begin        // N
                            x_32 = x_pixel - (368);
                            font_out = Nout_bitmap32[y_32][31-x_32];
                            font_in = Nin_bitmap32[y_32][31-x_32];
                        end
                        [402:433]: begin        // D
                            x_32 = x_pixel - (402);
                            font_out = Dout_bitmap32[y_32][31-x_32];
                            font_in = Din_bitmap32[y_32][31-x_32];
                        end
                    endcase
                end

                // BEST SCORE:    09
                else if (y_pixel >= 280 && y_pixel < 312) begin
                    y_32 = y_pixel - 280;
                        case (x_pixel) inside
                        [90:121]: begin        // B
                            x_32 = x_pixel - (90);
                            font_out = Bout_bitmap32[y_32][31-x_32];
                            White_in = Bin_bitmap32[y_32][31-x_32];
                                            end
                        [124:155]: begin        // E
                            x_32 = x_pixel - (124);
                            font_out = Eout_bitmap32[y_32][31-x_32];
                            White_in = Ein_bitmap32[y_32][31-x_32];
                        end
                        [158:189]: begin        // S
                            x_32 = x_pixel - (158);
                            font_out = Sout_bitmap32[y_32][31-x_32];
                            White_in = Sin_bitmap32[y_32][31-x_32];
                        end
                        [192:223]: begin        // T
                            x_32 = x_pixel - (192);
                            font_out = Tout_bitmap32[y_32][31-x_32];
                            White_in = Tin_bitmap32[y_32][31-x_32];
                        end
                        //space
                        [254:285]: begin        // S
                            x_32 = x_pixel - (254);
                            font_out = Sout_bitmap32[y_32][31-x_32];
                            White_in = Sin_bitmap32[y_32][31-x_32];
                        end
                        [288:319]: begin        // C
                            x_32 = x_pixel - (288);
                            font_out = Cout_bitmap32[y_32][31-x_32];
                            White_in = Cin_bitmap32[y_32][31-x_32];
                        end
                        [322:353]: begin        // O
                            x_32 = x_pixel - (322);
                            font_out = Oout_bitmap32[y_32][31-x_32];
                            White_in = Oin_bitmap32[y_32][31-x_32];
                        end
                        [356:387]: begin        // R
                            x_32 = x_pixel - (356);
                            font_out = Rout_bitmap32[y_32][31-x_32];
                            White_in = Rin_bitmap32[y_32][31-x_32];
                        end
                        [390:421]: begin        // E
                            x_32 = x_pixel - (390);
                            font_out = Eout_bitmap32[y_32][31-x_32];
                            White_in = Ein_bitmap32[y_32][31-x_32];
                        end
                        [424:455]: begin        // :
                            x_32 = x_pixel - (424);
                            font_out = co_bitmapout_32[y_32][31-x_32];
                            White_in = co_bitmapin_32[y_32][31-x_32];
                        end
                        //space
                        [460:491]: begin   // 0        
                        x_32 = x_pixel - (460);
                        if (score >= high_score) begin
                            case (score / 10)
                            4'd0: begin
                                font_out = zeroout_bitmap32[y_32][31-x_32];
                                White_in = zeroin_bitmap32[y_32][31-x_32];
                            end 
                            4'd1: begin
                                font_out = oneout_bitmap32[y_32][31-x_32];
                                White_in = onein_bitmap32[y_32][31-x_32];
                            end 
                            4'd2: begin
                                font_out = twoout_bitmap32[y_32][31-x_32];
                                White_in = twoin_bitmap32[y_32][31-x_32];
                            end 
                            4'd3: begin
                                font_out = threeout_bitmap32[y_32][31-x_32];
                                White_in = threein_bitmap32[y_32][31-x_32];
                            end 
                            4'd4: begin
                                font_out = fourout_bitmap32[y_32][31-x_32];
                                White_in = fourin_bitmap32[y_32][31-x_32];
                            end 
                            4'd5: begin
                                font_out = fiveout_bitmap32[y_32][31-x_32];
                                White_in = fivein_bitmap32[y_32][31-x_32];
                            end 
                            4'd6: begin
                                font_out = sixout_bitmap32[y_32][31-x_32];
                                White_in = sixin_bitmap32[y_32][31-x_32];
                            end 
                            4'd7: begin
                                font_out = sevenout_bitmap32[y_32][31-x_32];
                                White_in = sevenin_bitmap32[y_32][31-x_32];
                            end 
                            4'd8: begin
                                font_out = eightout_bitmap32[y_32][31-x_32];
                                White_in = eightin_bitmap32[y_32][31-x_32];
                            end 
                            4'd9: begin
                                font_out = nineout_bitmap32[y_32][31-x_32];
                                White_in = ninein_bitmap32[y_32][31-x_32];
                            end 
                            endcase
                        end else begin
                            case (high_score / 10)
                            4'd0: begin
                                font_out = zeroout_bitmap32[y_32][31-x_32];
                                White_in = zeroin_bitmap32[y_32][31-x_32];
                            end 
                            4'd1: begin
                                font_out = oneout_bitmap32[y_32][31-x_32];
                                White_in = onein_bitmap32[y_32][31-x_32];
                            end 
                            4'd2: begin
                                font_out = twoout_bitmap32[y_32][31-x_32];
                                White_in = twoin_bitmap32[y_32][31-x_32];
                            end 
                            4'd3: begin
                                font_out = threeout_bitmap32[y_32][31-x_32];
                                White_in = threein_bitmap32[y_32][31-x_32];
                            end 
                            4'd4: begin
                                font_out = fourout_bitmap32[y_32][31-x_32];
                                White_in = fourin_bitmap32[y_32][31-x_32];
                            end 
                            4'd5: begin
                                font_out = fiveout_bitmap32[y_32][31-x_32];
                                White_in = fivein_bitmap32[y_32][31-x_32];
                            end 
                            4'd6: begin
                                font_out = sixout_bitmap32[y_32][31-x_32];
                                White_in = sixin_bitmap32[y_32][31-x_32];
                            end 
                            4'd7: begin
                                font_out = sevenout_bitmap32[y_32][31-x_32];
                                White_in = sevenin_bitmap32[y_32][31-x_32];
                            end 
                            4'd8: begin
                                font_out = eightout_bitmap32[y_32][31-x_32];
                                White_in = eightin_bitmap32[y_32][31-x_32];
                            end 
                            4'd9: begin
                                font_out = nineout_bitmap32[y_32][31-x_32];
                                White_in = ninein_bitmap32[y_32][31-x_32];
                            end 
                            endcase
                        end
                        end
                        [494:525]:begin   // 0        
                        x_32 = x_pixel - (494);
                        if (score >= high_score) begin
                            case (score % 10)
                            4'd0: begin
                                font_out = zeroout_bitmap32[y_32][31-x_32];
                                White_in = zeroin_bitmap32[y_32][31-x_32];
                            end 
                            4'd1: begin
                                font_out = oneout_bitmap32[y_32][31-x_32];
                                White_in = onein_bitmap32[y_32][31-x_32];
                            end 
                            4'd2: begin
                                font_out = twoout_bitmap32[y_32][31-x_32];
                                White_in = twoin_bitmap32[y_32][31-x_32];
                            end 
                            4'd3: begin
                                font_out = threeout_bitmap32[y_32][31-x_32];
                                White_in = threein_bitmap32[y_32][31-x_32];
                            end 
                            4'd4: begin
                                font_out = fourout_bitmap32[y_32][31-x_32];
                                White_in = fourin_bitmap32[y_32][31-x_32];
                            end 
                            4'd5: begin
                                font_out = fiveout_bitmap32[y_32][31-x_32];
                                White_in = fivein_bitmap32[y_32][31-x_32];
                            end 
                            4'd6: begin
                                font_out = sixout_bitmap32[y_32][31-x_32];
                                White_in = sixin_bitmap32[y_32][31-x_32];
                            end 
                            4'd7: begin
                                font_out = sevenout_bitmap32[y_32][31-x_32];
                                White_in = sevenin_bitmap32[y_32][31-x_32];
                            end 
                            4'd8: begin
                                font_out = eightout_bitmap32[y_32][31-x_32];
                                White_in = eightin_bitmap32[y_32][31-x_32];
                            end 
                            4'd9: begin
                                font_out = nineout_bitmap32[y_32][31-x_32];
                                White_in = ninein_bitmap32[y_32][31-x_32];
                            end 
                            endcase
                        end else begin
                            case (high_score % 10)
                            4'd0: begin
                                font_out = zeroout_bitmap32[y_32][31-x_32];
                                White_in = zeroin_bitmap32[y_32][31-x_32];
                            end 
                            4'd1: begin
                                font_out = oneout_bitmap32[y_32][31-x_32];
                                White_in = onein_bitmap32[y_32][31-x_32];
                            end 
                            4'd2: begin
                                font_out = twoout_bitmap32[y_32][31-x_32];
                                White_in = twoin_bitmap32[y_32][31-x_32];
                            end 
                            4'd3: begin
                                font_out = threeout_bitmap32[y_32][31-x_32];
                                White_in = threein_bitmap32[y_32][31-x_32];
                            end 
                            4'd4: begin
                                font_out = fourout_bitmap32[y_32][31-x_32];
                                White_in = fourin_bitmap32[y_32][31-x_32];
                            end 
                            4'd5: begin
                                font_out = fiveout_bitmap32[y_32][31-x_32];
                                White_in = fivein_bitmap32[y_32][31-x_32];
                            end 
                            4'd6: begin
                                font_out = sixout_bitmap32[y_32][31-x_32];
                                White_in = sixin_bitmap32[y_32][31-x_32];
                            end 
                            4'd7: begin
                                font_out = sevenout_bitmap32[y_32][31-x_32];
                                White_in = sevenin_bitmap32[y_32][31-x_32];
                            end 
                            4'd8: begin
                                font_out = eightout_bitmap32[y_32][31-x_32];
                                White_in = eightin_bitmap32[y_32][31-x_32];
                            end 
                            4'd9: begin
                                font_out = nineout_bitmap32[y_32][31-x_32];
                                White_in = ninein_bitmap32[y_32][31-x_32];
                            end 
                            endcase
                        end
                    end
                    endcase
                end

                //   MY SCORE:    03
                else if (y_pixel >= 350 && y_pixel < 382) begin
                    y_32 = y_pixel - 350;
                        case (x_pixel) inside
                        [158:189]: begin        // M
                            x_32 = x_pixel - (158);
                            font_out = Mout_bitmap32[y_32][31-x_32];
                            White_in = Min_bitmap32[y_32][31-x_32];
                        end
                        [192:223]: begin        // Y
                            x_32 = x_pixel - (192);
                            font_out = Yout_bitmap32[y_32][31-x_32];
                            White_in = Yin_bitmap32[y_32][31-x_32];
                        end
                        //space
                        [254:285]: begin        // S
                            x_32 = x_pixel - (254);
                            font_out = Sout_bitmap32[y_32][31-x_32];
                            White_in = Sin_bitmap32[y_32][31-x_32];
                        end
                        [288:319]: begin        // C
                            x_32 = x_pixel - (288);
                            font_out = Cout_bitmap32[y_32][31-x_32];
                            White_in = Cin_bitmap32[y_32][31-x_32];
                        end
                        [322:353]: begin        // O
                            x_32 = x_pixel - (322);
                            font_out = Oout_bitmap32[y_32][31-x_32];
                            White_in = Oin_bitmap32[y_32][31-x_32];
                        end
                        [356:387]: begin        // R
                            x_32 = x_pixel - (356);
                            font_out = Rout_bitmap32[y_32][31-x_32];
                            White_in = Rin_bitmap32[y_32][31-x_32];
                        end
                        [390:421]: begin        // E
                            x_32 = x_pixel - (390);
                            font_out = Eout_bitmap32[y_32][31-x_32];
                            White_in = Ein_bitmap32[y_32][31-x_32];
                        end
                        [424:455]: begin        // :
                            x_32 = x_pixel - (424);
                            font_out = co_bitmapout_32[y_32][31-x_32];
                            White_in = co_bitmapin_32[y_32][31-x_32];
                        end
                        //space
                        [460:491]: begin   // 0        
                        x_32 = x_pixel - (460);
                        case (score / 10)
                        4'd0: begin
                            font_out = zeroout_bitmap32[y_32][31-x_32];
                            White_in = zeroin_bitmap32[y_32][31-x_32];
                        end 
                        4'd1: begin
                            font_out = oneout_bitmap32[y_32][31-x_32];
                            White_in = onein_bitmap32[y_32][31-x_32];
                        end 
                        4'd2: begin
                            font_out = twoout_bitmap32[y_32][31-x_32];
                            White_in = twoin_bitmap32[y_32][31-x_32];
                        end 
                        4'd3: begin
                            font_out = threeout_bitmap32[y_32][31-x_32];
                            White_in = threein_bitmap32[y_32][31-x_32];
                        end 
                        4'd4: begin
                            font_out = fourout_bitmap32[y_32][31-x_32];
                            White_in = fourin_bitmap32[y_32][31-x_32];
                        end 
                        4'd5: begin
                            font_out = fiveout_bitmap32[y_32][31-x_32];
                            White_in = fivein_bitmap32[y_32][31-x_32];
                        end 
                        4'd6: begin
                            font_out = sixout_bitmap32[y_32][31-x_32];
                            White_in = sixin_bitmap32[y_32][31-x_32];
                        end 
                        4'd7: begin
                            font_out = sevenout_bitmap32[y_32][31-x_32];
                            White_in = sevenin_bitmap32[y_32][31-x_32];
                        end 
                        4'd8: begin
                            font_out = eightout_bitmap32[y_32][31-x_32];
                            White_in = eightin_bitmap32[y_32][31-x_32];
                        end 
                        4'd9: begin
                            font_out = nineout_bitmap32[y_32][31-x_32];
                            White_in = ninein_bitmap32[y_32][31-x_32];
                        end 
                        endcase
                        end
                        [494:525]:begin   // 0        
                        x_32 = x_pixel - (494);
                        case (score % 10)
                        4'd0: begin
                            font_out = zeroout_bitmap32[y_32][31-x_32];
                            White_in = zeroin_bitmap32[y_32][31-x_32];
                        end 
                        4'd1: begin
                            font_out = oneout_bitmap32[y_32][31-x_32];
                            White_in = onein_bitmap32[y_32][31-x_32];
                        end 
                        4'd2: begin
                            font_out = twoout_bitmap32[y_32][31-x_32];
                            White_in = twoin_bitmap32[y_32][31-x_32];
                        end 
                        4'd3: begin
                            font_out = threeout_bitmap32[y_32][31-x_32];
                            White_in = threein_bitmap32[y_32][31-x_32];
                        end 
                        4'd4: begin
                            font_out = fourout_bitmap32[y_32][31-x_32];
                            White_in = fourin_bitmap32[y_32][31-x_32];
                        end 
                        4'd5: begin
                            font_out = fiveout_bitmap32[y_32][31-x_32];
                            White_in = fivein_bitmap32[y_32][31-x_32];
                        end 
                        4'd6: begin
                            font_out = sixout_bitmap32[y_32][31-x_32];
                            White_in = sixin_bitmap32[y_32][31-x_32];
                        end 
                        4'd7: begin
                            font_out = sevenout_bitmap32[y_32][31-x_32];
                            White_in = sevenin_bitmap32[y_32][31-x_32];
                        end 
                        4'd8: begin
                            font_out = eightout_bitmap32[y_32][31-x_32];
                            White_in = eightin_bitmap32[y_32][31-x_32];
                        end 
                        4'd9: begin
                            font_out = nineout_bitmap32[y_32][31-x_32];
                            White_in = ninein_bitmap32[y_32][31-x_32];
                        end 
                        endcase
                    end
                    endcase
                end
                
                // NEW HIGH SCORE!
                else if (y_pixel >= 180 && y_pixel < 212 ) begin 
                    if (score > high_score) begin
                        y_32 = y_pixel - 180;
                        case (x_pixel) inside
                        [40:71] : begin                  
                            x_32 = x_pixel - (40);
                            font_out = Nout_bitmap32[y_32][31-x_32];
                            countcolor_in = Nin_bitmap32[y_32][31-x_32];
                        end
                        [74:105] : begin                  
                            x_32 = x_pixel - (74);
                            font_out = Eout_bitmap32[y_32][31-x_32];
                            countcolor_in =  Ein_bitmap32[y_32][31-x_32];
                        end
                        [108:139] : begin                  
                            x_32 = x_pixel - (108);
                            font_out = Wout_bitmap32[y_32][31-x_32];
                            countcolor_in =  Win_bitmap32[y_32][31-x_32];
                        end
                        //space
                        [170:201] : begin                  
                            x_32 = x_pixel - (170);
                            font_out = Hout_bitmap32[y_32][31-x_32];
                            countcolor_in =  Hin_bitmap32[y_32][31-x_32];
                        end
                        [204:235] : begin                  
                            x_32 = x_pixel - (204);
                            font_out = Iout_bitmap32[y_32][31-x_32];
                            countcolor_in =  Iin_bitmap32[y_32][31-x_32];
                        end
                        [238:269] : begin                  
                            x_32 = x_pixel - (238);
                            font_out = Gout_bitmap32[y_32][31-x_32];
                            countcolor_in =  Gin_bitmap32[y_32][31-x_32];
                        end
                        [272:303] : begin                  
                            x_32 = x_pixel - (272);
                            font_out = Hout_bitmap32[y_32][31-x_32];
                            countcolor_in =  Hin_bitmap32[y_32][31-x_32];
                        end
                        //space
                        [334:365] : begin                  
                            x_32 = x_pixel - (334);
                            font_out = Sout_bitmap32[y_32][31-x_32];
                            countcolor_in =  Sin_bitmap32[y_32][31-x_32];
                        end
                        [368:399] : begin                  
                            x_32 = x_pixel - (368);
                            font_out = Cout_bitmap32[y_32][31-x_32];
                            countcolor_in =  Cin_bitmap32[y_32][31-x_32];
                        end
                        [402:433] : begin                  
                            x_32 = x_pixel - (402);
                            font_out = Oout_bitmap32[y_32][31-x_32];
                            countcolor_in =  Oin_bitmap32[y_32][31-x_32];
                        end
                        [436:467] : begin                  
                            x_32 = x_pixel - (436);
                            font_out = Rout_bitmap32[y_32][31-x_32];
                            countcolor_in =  Rin_bitmap32[y_32][31-x_32];
                        end
                        [470:501] : begin                  
                            x_32 = x_pixel - (470);
                            font_out = Eout_bitmap32[y_32][31-x_32];
                            countcolor_in =  Ein_bitmap32[y_32][31-x_32];
                        end
                        [504:535] : begin                  
                            x_32 = x_pixel - (504);
                            font_out = ex_bitmapout_32[y_32][31-x_32];
                            countcolor_in =  ex_bitmapin_32[y_32][31-x_32];
                        end
                        endcase
                    end
                end

                // 카운트다운을 위한 카운터
                if (clk_counter_end == 25_000_000 - 1) begin
                    clk_counter_end_next = 0;  // 카운터 초기화
                    if (countdown_end > 0) begin
                        countdown_end_next = countdown_end - 1;  // 카운트다운 감소
                    end else begin
                        if (score > high_score) begin
                            high_score_next = score;
                        end
                        state_next = IDLE;
                    end
                end else begin
                    clk_counter_end_next = clk_counter_end + 1;  // 카운터 증가
                end

            end

        endcase

        // 일반 디스플레이는 검정색 폰트, Win은 Blue, Lose는 Red
        ////////////////  WIN  /////////////////////////////
        if (w_mid & ~w_in) begin
            red_port   = 4'h2;  // Red
            green_port = 4'h9;  // Green
            blue_port  = 4'hC;  // Blue
        end
        else if (w_in) begin
            red_port   = 4'h6;  // Red
            green_port = 4'hC;  // Green
            blue_port  = 4'hF;  // Blue
        end 
        else if (w_out & ~w_mid) begin
            red_port   = 4'h0;  // Red
            green_port = 4'h0;  // Green
            blue_port  = 4'h0;  // Blue
        end


        ////////////// LOSE //////////////////////
        if (L_mid & ~L_in) begin
            red_port   = 4'h8;  // Red
            green_port = 4'h8;  // Green
            blue_port  = 4'h8;  // Blue
        end
        else if (L_in) begin
            red_port   = 4'hF;  // Red
            green_port = 4'hF;  // Green
            blue_port  = 4'hF;  // Blue
        end 
        else if (L_out & ~L_mid) begin
            red_port   = 4'h0;  // Red
            green_port = 4'h0;  // Green
            blue_port  = 4'h0;  // Blue
        end


        ////////// 32 * 32 알파벳 & 숫자 //////////
        if (font_out & ~font_in) begin  // 테두리 검정색
            red_port   = 4'h0;  // Red
            green_port = 4'h0;  // Green
            blue_port  = 4'h0;  // Blue
        end
        else if (font_in) begin
            red_port   = 4'hF;  // Red
            green_port = 4'hD;  // Green
            blue_port  = 4'h1;  // Blue
        end 
        else if (R_in) begin
            red_port   = 4'hF;  // Red
            green_port = 4'h0;  // Green
            blue_port  = 4'h0;  // Blue
        end
        else if (Y_in) begin
            red_port   = 4'hF;  // Red
            green_port = 4'hF;  // Green
            blue_port  = 4'h0;  // Blue
        end
        else if (B_in) begin
            red_port   = 4'h0;  // Red
            green_port = 4'h0;  // Green
            blue_port  = 4'hF;  // Blue
        end
        else if (countcolor_in) begin
            red_port   = 4'hE;  // Red
            green_port = 4'h3;  // Green
            blue_port  = 4'h3;  // Blue
        end
        else if (P_in) begin
            red_port   = 4'hF;  // Red
            green_port = 4'h0;  // Green
            blue_port  = 4'hF;  // Blue
        end
        else if (G_in) begin
            red_port   = 4'h0;  // Red
            green_port = 4'hF;  // Green
            blue_port  = 4'hF;  // Blue
        end 
        else if (White_in) begin
            red_port   = 4'hF;  // Red
            green_port = 4'hF;  // Green
            blue_port  = 4'hF;  // Blue
        end
        


        if (cha_1 & ~cha_2) begin
            red_port   = 4'h0;  // Red
            green_port = 4'h0;  // Green
            blue_port  = 4'h0;  // Blue
        end
        else if (cha_2) begin
            red_port   = 4'hf;  // Red
            green_port = 4'hf;  // Green
            blue_port  = 4'hf;  // Blue
        end 
        else if (cha_3) begin
            red_port   = 4'ha;  // Red
            green_port = 4'hf;  // Green
            blue_port  = 4'h7;  // Blue
        end 
        else if (cha_4) begin
            red_port   = 4'h6;  // Red
            green_port = 4'h9;  // Green
            blue_port  = 4'h6;  // Blue
        end
        else if (cha_5) begin
            red_port   = 4'hf;  // Red
            green_port = 4'hc;  // Green
            blue_port  = 4'ha;  // Blue
        end
        else if (cha_6) begin
            red_port   = 4'hf;  // Red
            green_port = 4'h9;  // Green
            blue_port  = 4'hb;  // Blue
        end
        else if (cha_7) begin
            red_port   = 4'hf;  // Red
            green_port = 4'hd;  // Green
            blue_port  = 4'h3;  // Blue
        end
    end

endmodule